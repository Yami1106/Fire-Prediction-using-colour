PK   6f�Xn�
�$  ��    cirkitFile.json�]]��6��+]��n��� 	�[��Ԧjg��l�>�.?��iK=ju����}AR����=t��+�������.>?/v�/�fUlw��j���nw2Z.>d��Sv�[�\<�7��v��]��aq���9���P����|k�YE���ˠQ�4-�<�d��*�
S�,)Vb%wo�/�G�l��l\�Rl\�
��b���b�9p�*fs�"�U���E+���E��́�`c?P�!,@���J��l˂.��?`�!,~�dCX��Ɇ�,�a�aY�'²��N6�[�c'²��N6�eh�c���N6�e���l˂;��?v�!,~�dCX��Ɇ�,��Ӂx�~�v�.[ߓ�����>ۭ��ٛ�p��/L8�{+���j�_�Y�Wu�qeK� �Q�R���C)B���1�?��8�f�X�C�I,;��`m������.��� �z�*Ě=Ě�Nbى���Ncme'���*��.���NbىU��]����Ĳ�k�k;(;�e'Vk;����Ĳ�k�k;(;�e�̢����|�O��5��`��tfNM$87����O��5k.`���,?	�׬���4��$�_���8���`~�
�~���O��5k�`���,?	�׬����<��� ����R��2�J��6ub��$�UZ�4V��b����-��`�I0�f<�N]\~����eR�UE�t^6`����42O�B0]M��Y����`��~W7%oY�ٮ 6=z5��N�8aR��	�O�rݤP�uT��m=60�6Ah�H��K�D|��Z
�ka�I0�f_�~�\�O��5;z���ZX~ً̯�8���`~�.*���������Hq��%"ε8�r�]�K�s�ц�d���\g�,�
tf��TE�*�R�(5}*���f�IT$�JoƠ��i<���ቷ���N���)w��1g3Wȱz©Yqj�x{��T��o�z{������'�z?���#<W�OɊY���S���<���Qg:�s@fj�ez�s(e��L�o�\=A�
��鏩�3�������g%���t]�|��n����g�)�TM�.gZAP����^&IiT!�F{*_T!����_�cP�yu©Zq]�P�:�2�Mu���<ȳ���Q��u�E�k���aé�gR�)�fũY�RaRվW�V�o,F�Z���9U��δ�}��jV�)Y�J5%���j_�K�:eU��\h��l�ȩ�μ�$Zݬ��{lV@�=5+���w2�T�/�O22����T1�	idN��c��X��I�\����L��}�O��}�95`0����Ԁ���כ���}�9q�ω.���8��T��ʉ#|NվPF�q���2⨏S5/��<�ەSG}��Y�ͼk�|�S5+��:MɊg����J��v%�K�����펯O��F���$
��c�0�S�F �v�����b��Z�[#P�y�ajp1�@@�.��U��0uZ����ڸ����QH��.�,vKX�F!u�� N��-a�ԩ�8�b��qR�����
�QH��/�n����⸂�qR�����
�QH�0�,�+XG!u:� N�8�`q܇��mO{�QۃTWQx��?@Qa\]�`8*Юspu��1�醣�:WWUx�4��i��g�1v���X`��l0����pT�]���J
c,�?�G�u���0����pT�]���Jc,�?G�u��L1����pT�]���Jc,�?G�u���1h?O��	���s��>a��k��k��k���Q��"m;O�5��d<,Ҷ�_��PU��"m;O
6��e<,Ҷ�a��Pc��"m;O*6��f<,Ҷ�c��Pq��"m;OJ6�1G�� �l;OV6��f�
�<y�#wZ�g)l��xX�m����"b�#r��L+b3-�͓�9�xX�m����B�v���:a��l���xX�m���fa;�܌�E�v��l���xX�m���fa;����E��e�γV�H&�a��u�Bl�u�	Ӆ���M�Lp�쾞�z@��p���@iw'�N�b����r�ȳSw�R1 �w<�
�b�}}綮3F�<8)����Lq�UIŁ�8��������\�J�����ZZs`0^�;r��0�s�
�a�E/�j�� �2��ц�<>�����?U�wܺT9�񷉪�{ቈ���1��o;�FTiچ��ӂ��>QTg��<U2v�M]�����c�a�@��Dg!���il��0Pڠ����<�W�R��,���.dʺ�9-�F̺2)�w�ѫ}����R�UE-Ln�M�67й�����Eu]rZ[8�YՍ^�D�>�P5��&Us<�Q�,ǳ8�(�xFI�w�V��Pe�����s�W�
+��Jd���n�,x8�/���0Y�p<�E�#0Yp<����;m�l�x�M����rz��6Yo|MV�{�y�{�g�
 ����������uBy �.�0u���˫ �@@�P��ʃ0uByF �N(��	�A��:�<#�A("qQ�aq[�7
� ������QH�<'X��� �B:�a8�b��q�A(�	�,���ByN��7n ��
�QH�<'XW�8�B:�a8�⸂�q�A(�	�,��� Byh�n� u@(�
�: ��F�u�By8'mШ@���u@(b�h�9��A,���A��:��<���5hT�]��: ���s��
��\�� pNՠQ�v���P�Ή4*ЮspʃX�9M�F�u�By��<	�+=��ϓr��vH(���Li�<y�+=�E�v��k�CBypX�m�I�fa;$��E�v�l�CBypX�m�I�fa;$��E�v�Tl�CBypX�m�I�fa;$��E�v��l�CBypX�m�I�fa;$��E�,̓���vH(���<y�,l����H�δ$6O^�J��a���'/���Pi�y�Y�	��a���'/���Pi�y�Y�	��a���'/���Pi�y�Y�	��a���'/#��B(�����}�Pų_�
�<>�gO�By|Ͼ�+���(�����`0��;v�P ����Q��`0>�;6t�P �a��w���< Ƌ}M���`��w��< �E/&��Q.�0Y(����r�u"卣P���(��B�E!��Q.>Y(��r���By|��Q�,��G�3�By|���.���x���+]( �q�ˣW�P�b;����([�,��G����(C��\�2d�<�ׁ�㽗�]( �q`P���#Ӆ� 0'��#Ӆ� 0�^�ei���~Ulﷻպ�uq����zW=�*W��j�+�����[Ƅ���|b#r�<ԁ.��r� s[wQ�$��C������A*���EEG8*����Ľm*��k^�8�x�ꉎ�:γT�
ҬI�A�+�JV�֡0��Z���C���]d�����C���Qn�΋s��x��~ʡ��9Us���"_�:5a�RTih�(%k[uUY��<�JQ&f����j�۽�S�=�T����D��9<�I�[U�;�z��)g\���m��ѧ�T�
���P�9����U+O8$� p�8�C��p ��4G�p�_�UhK^<*�a*q݌G�6x'.x�������۷8����'9n��S�"�f����w8G�:�,���d,�5DV՞~���Ȫ��Y/V�OxUs>LexUs�Ɩ��|.��˪�3 �.�r�f=6/�����8�L��'�Ɉ;t��8��#pG���qK4g�S�������W�v���/U��6��j�[�������g�m�ѫ���������^wk����GNt�]�G�#�L�(�WY��3B�[Z��|ɷ	w�� ���g�]��3�.m�c�뼺cQ�u^]6#v��_]6O�M^�3�6#v�0�*��6�:�#l��(�p�o}�m|B��L�d�"1�o���ʻ90���:^1�]�k���s1eL6�e�;�:ܱ	����W
6lJ��I6#��{�k�y������߯8a��f-q�(ܽ��V�V?���&,�m�|�ݟ��^e(�O�{A�m�[B���;C�~�� :���>�Q}��|�]�|�ͣ �=� ̭� �� ̍� ��� �m� �ݦ �M� 
ܽ�|
�-�|ܝ�|��|�}��r{*�$�]��܀�Y�O��g�2Xd��i�ٮ�پZ�=����}�߮������K]����|k�R����)ݩ��i?2Y�!:�H&6D�=�d�����B�ZeLl�j�1Y�!D���d�����B�ZmLl�i�q�"z"�' ~J@ �c�N���C% ��1D'�����H������ �R	�|щry ��S>��d�<�QĀO ��1D�u.@<U�x�����< �T�)Ct_h�� �S��.���m9_���u��b�9�Xwq�G�0x ]�M���|=�iN,?	�'V·rqx�a�9��{'��w���4��Q\��c�I0?�r��Ã��O�����[�~X~�O������ ���`~b�|�������	H<����$��X9ߜ��A��'����s�x���J4�f�mCxR�J�i�D�%���J4�f�mCt6f(���"��	��D3lV��6Dg%`�ͰY�C����J4�f�mCtvf(���������ϧ�aZ ��Ht�f(��sN
��Ǿ��"��*`���Ƥ�,��=[�sq@�[�-��tR��IM��)���I�˰�>���I�9��D3lv��m��q�%�a�smCt�f(���{06D�8`��P8�P@������u>Ƥ��/�7�ðgR��������P3Q�d��d��!�T�~�L����l.�x��)t��Gg���=����gk����-�S���>]6�	�uP�X�T ���Az�,K��ـ<]1�!���q��=
15�q��=|0���v�^��T͹n���pv�O�:���|��u,AգF� ��L�d���I��p#oQY��B���&+�Qc0Qon<Ϙ,�ՇcIL��ҋr�%��:
K�G�p��pG,iw���r�,,��q$�R������Z����}1�Ő�����

9x,�&��P�w���3~�d�V����:7�ܒ��C�|�b[T�#*gQ=�(�Eu<������'��(��-U\���R�"��-U���iP����U���kP����U8�:`��`RG,TQKꐅ*QI��������|��\�ܸ.�2���ȕQ�����E�V�+4�g�J5�ؘ�1W��kѸr^ڠо���׶y�P�u[���Q���Ƕnֆ�6�!�|m����m��O�/(�i{%�s�����!��ho��0P6��Q<��4�{�hO�m�}�^+[��(z:�IO�4��F��05�6�Æ���	9l���;�a�*:����WLv}M}�]��k��;�;�־��p����K���׬9s�;��_C��!��_C��!��_E��a��_E��a��_E��a��_E��a��_E��a��_E��a��_E��a���0���l+����a�b�7:�h��>�Æ���
pذ�1��V4�~C�a3G_��	8�X��m��/V��8d|��k|s�ee_��_�gyu�L��ޟ���O���i��y�$�K�pI���åн���{):\��K��R�^J���9\2��p)u.ɣ5�k�l��h�D"]�ȣE�ky4�tm"�6��Q��(ҵ�<ZE�f�G�H�.�h��E�\��g?q�vQ�]��.ʵ�:�E�vQG�(�.�h��E�\���]�?�;��߯N�?כz��_?�۹Q��vc�)��s�T������xD"Y����ofUs!�ȂDT&С���e �04�v$i�5�������ZR���􏶿KU����n��(2*�6�"�q]Y�����;,d3�O�UY8��?=�Ӷ�	E��myi�� K�*E,eQ|F.��*}6-)���h81-������*���9�>�>�g�s��7��C�ۯ�f��z��`���vcH-o�$�{</��n�	�~e����ci�J�i����MC�AZ�:�tb�Z�y�-N����=�5��b�y�g��"-�,��ڢd�Ek�b�+����md�$��XF�mb[W��O����NΊ�d�X�HŒ�.�*R1���r���)��S�)]|ԦT�\��)d.��v���UM���s�����4X�m��bn;h��r�v�sj���T���.�4�p����-7��J|D)�>��+?T���@����Zʵ1�l���jYo��j���n��>V�w����Ňw��źl��8��Ў��<t�� e��a�a��m��ׇ���������ݽ�$u�i D��1��ܘ8�3��\k%M����r_��0-�0��M��A�JFi)D%L�|ߏ������U���3;H�U�H��	�2�-DR�����{��7�Q5�6���M�z�$�Xߗ'��7�\Z�(��ȳ�h�;XxQI�a֙)��v�����js����3����*��� ��PV�LE��(��o�S6�(E�W����J��2I��Y�3�F���ï٦�����_��;|*����o��ElK�^���-��~y���/o���?��\m��[�lw�o�rW=>�,�R+����Հ��ڛN]M�2ODm;�B��^m�ΤUn��B&�(�*�|��:7y(�266��Tl�]q"���C�䃮f�aa��V'�@�ydQ-SV�.L����ZG"/j�ՙ�BVA������u��:���Պ��w�_�����?=�˿�|~�nss�����n~�>�+7M�ծZ��7����֎W�li�ߗ��~�����70����Uy��)X����*����e)��.��{�������I�e��P��v�������S��>���6���	6�_�(ϖ|��֛f��������\���?5?�$lҭ��ڎX�_���~�|oA�f_<=V�?���}���]�����*�O���m���?YG�����oˬ�=��7?nʧ����|plS m�%ɡc���=B;65�����q�K�ihG�M~r]�P���eX�Q�����Շ0<¦�Z���}X`��[�_Y����׸L/�P�6�Q��e�����q�;��S�$0��k����Z��<uT6���ԒK) mm"��-)�y&�r�k��}��>��m�� �X�֤,�T�FF"���Y�J�6�ֶ#3ebS-�4AlL�ʄ�fsʮ0�SJ���\���6��WS}��+�Ne���(h�?I���֎J��׶I��;Je�n�:Z�La�Qe���*�;b��GF$J;Z?��vR&l�O=C[oѽ��݇M
(�0�~���rZ�}#i�8B�9��D@CL{��)IE+��x��&QD�K���р�!U.���˟�r��o{�&ڗ��*��>cSQ��&J����J��Q`3�"���,ȴLd3��"Ez�H[k��_���|�j ���:C7���ȹnN�7Ǎ�������Dh�I�Xe�Ǥm�g up��\"^�l�\��XK��un!mrԕK<����H:>�M���mlj����ib�c◑�p�68Eփn�-���m��`��g�f����4����[���L�ͬۧ�fo�c�T���}��#�xK�] ���m�L���ꚾ��~�BaG��U�����QW�DCF�~�}ڔ�e��}��ٛX�Mv�.���i�&�DM��i]�?4JۗIǺ�凪]��[�6�����o��͡���P��=�a��U��o^W���#����M�}�ݵ��7B$e�M��(�ۿYo���ỉ�M9�E��B�O?C�Y�?��=lכ��l������ݻE�h�S����s;^|l~{����ٔ��|����t�qt����Fr�H���n���S�5�*�����\�vR�	�5&Л���>��J��ٵz��O-�����Q(S�5�;TH����w���tzS��l9gu\Y�9�y�@�z;"^�Vʦ~$����:�5Ĉg���]E�{
��D�9[��x�y}��/�B���T8���Ta��\�6�"�f��D�i���� `��p������&=�j15\��bN�a�����i��b���C��Н�b�Ч����G�i�{9�Q�t��ڨC�t��S�9"�0�X�H1P+h�@��!���"c��5��1z�-^8�nA:~u��i\�(/��N��k��~ᤰ��r�H�3�r נW�-���Δ�\���e"�-�/f����1��h�ES��{hg�I�)���tg�@�0�2��Ԝ�l�g�[�yI��^0 ӴV����IV� ��'̱N��j���Xϗ�V�բ���k�Ljc]��˂4��9�Z��D:��Q�j4��C^�A��75=[����Sl��u?E!#�Gl�2̡�1��L�@�ǅ��*zS��<oF��S����|�X�=��P��q���C�C_��;ƣG����Äҹ8ň�a�0Ye��A[ޥ�ʠ݃��;��T�x��2��b�v��k�Q���u����Gb�{`��*�8nv:���=��<�ӢG��=�$J4uڜ���s����%��=����G�~1O�Z��#���u]C�Z9��;U	�o��7�=�7���G����SZ��/F�V&%/���p݃�yh���q�x�=�b�����N1�{�e�ԽeDq8�z2Tj�ȫ�C�w���чS���?�bTɛ�� �]�D�>����-O�7�A����G�~1O�k�̩S�� I�u.�� �Sp��j���Pϸ{�y�=�ŏ~1j��u	Mn��=s
�W͜���w�~1O�'��G�y�4���p�T�gN�����#|F�b�v7����sIt�} 'N%z�;q*��9}>�������_z1b�O�*J؍�;W�=w�+vp���'�O�;��b1M�O����C�G]�9lU��0�ް��5|� <;E.z������<}N�C����I}M���-���	�xG1=���r��U��T�\8����1�)��]h=�B�����C�L`7��D}�s^�l���1����
��9���뼧�1X���T�1�W�uv���k��a�?U��l�������؈�}�8��n��U��}�X����ŗ�PK   6f�XG�~��  � /   images/0739a1b1-a163-452a-a325-ab452d55b136.png�y8�m?�r�J�M!*IY��Ie�^Y&������[�d�cb�0��d�1̒,�ٲ�L������������|�|�4}��>�r}��|��mn$�_l��mۄ�o^�ܶM�i۶]&{w-�����A���{����� ��n�m�&�I����em4�6�l����
�*y�����x(����WŶm;����5��9t4Gb&��Ȳѹ�}��OܜΉSٱ������b��MT�}�L�1HƸD���?j��i͘�ǰf�	�A��{�ξ�[_����J�z���r���٢w��/5a��t�I��ե�EnhǶ-?����'m�ں-��Ǔ[�n�-��v<����xN��J�h���e3��2������7��=V��)u!";G?�� ��<�|K0�yY���I2,���^)�Ϭ���Ev�p�����������d���4���dK;!-�L�^�$Cx�䐦W��k��E���9謗	* P��ϕ�����S�����0C���~�?��$Ǖ���φ%mXJ����{���w/�y|
�T!��;��G����쳄�[�����⩧�U�6}3���6��{�[$��ab1�P��~z�3������Y�q(�V�f��¦�&	�� ��l.Z��s9�2SH�W�ơP6�[��SnT�QokF!s�Ǔ`��� 6rl�������fI�:�v�K�|l��%����)�m����}gw0�6=y�dk��?�/������<�w�}l��جJ���s�+����������6����Í�͍{3�����"R-33�	a\yoU+����̡-�߶~�S���v�ѯ�f��nY7�߼�K�pE߬�����f�J�\t���+"D�,�����AGf�H��X��i���&���oց���A{10�^���l����UL&0���ٵ?���E�)�Q�5��s�=[�,�8�v�Y����>\��>\+sS�N��88y��</�!-Ot�HS�/'9��q�ZwuR��
���ӝ�v�����xS>edf5�Ի`��Z��/�j�3�QM�/
�1Q �wH����G�h�p���"[�|���fi�h.��-
��f�:�[<?>gh8)�2d����q���j�GZl��Ϩ�4.{��F���Hq���5�1͸�m2�2~�l����]I���J�&k�-�x�T�/�O�z�5�k����8��JdX��a9�<��V��\�����R��9�����0�TƦ%r�hm�[o���b�Pԓ��YپQ5Y�� �>[Զ�f�UG~����bhA�A	���6��,-��:[��Y����p���m���k���A��p�ʂ�K��&�{sdJ;?=3�O�	}�Ij�>>wE�Ws20NJ]=X�uq�g�j����bN���|�G����Q�s˪�r���W��ӕ������7�[����v�ЂF�K^��FY�{��s��ʻ��R�:i��D{��x�����T�Dr��j�M�s3�����:u˙��[�.�[Im}�v8��0��d�Y�S�ܷ�BW�V�F��V�E��V�
���355;����҈�RW&/�+�'��]W�e����v�@$�Y��=�Vܲܽ��ٳ�6�tinb��[s!ޞ�C����<_��iG�Gn���_a+*�� ]>��-u��{\lrǹ��x�|�b�ߕ��?e��@�㕸�����[�`J�p-��i��m�'���n��:l�xm�pd�l�em,W0Q�:��"�A�fXDyP��pOTG^uPiN��c��+l����~ŭdyώ�ȂrZ�����?���A�Xc|O���/�Pc���>���tx/��g�N8^xai=���
\�ΟNXi��@�l��]Q�0��!a�+ץ���q�����`Vq,�o"�B8a�i���Itq�����1C�06�J��J���
�<-VTy�����kQ
�ɍ������p�F����Ϝ����r�}��O��u�~�Ar�u�����Wc~2�ƪ����@�m�����
&�H�;7��.2g�>)l!�(�|�v�z��[�TJ�й��#�J�:F���R���:oȼ�>33�w��vå"����P|�?{�&��#�H��+���#��<o��Jڐ(-�������&�Mt^��R��|٢����q`�g��c��j��02���)����F�;W������+�xR��:P��/�ސc�H���\k�Ý�/���d�����^� u �Ƚ���c��������-6yK�.�d�j��܉�x�������7�.{��"�'�>����K�۰o�g����m%���UY�> �/��
zo��X{_�v��Kû��q��Ŧ�ү2#G�_Z&�k3��x��r��2#zל���@�[��װ��^_�L�#/=lql�X4Xm������nq�p�7ME]�A��J60��e��ogU.Ė�FՄ�W_Ћ�[cT���l�hze< &��x����/{�"�Lv��
��= з$:��Ln�_�|_�!��ɬK{U���G��Jak�6����������R3Ć��S�ۿE$��|��ӝ1��E}��q[s<w�R��.�$����V�P���Lկ�0e�YK�9��qO_L���p��Tu��/8�ˊ��Z��]��A�@(�^�1���s�z��'�l��x�}u��A���<�� m������j��1õ��B��iB��	�A&q��6�t���+�cQ"M	��յN�I/&�'9�˹��Vv�t�R��FAD�/��"������N��+�',��Z.����xT�;(a��C��?����Drɴ��J@a��m�e��h?-����b	���M8=�^����=�ӽ�b/��Y:#�3���rp`��$G7��0_��s�N���vo���B��
]\�R�	�e�1cٝ)z)A���۹����E;DO�V$���t+˾C��@;�sA����.���8yQ\��Gwz�O/9s>u��ř����e�5o��e=���qפkx�t������]�o�O��V��f(�\z/�x�@P�p8��R��fU�j�nL�`v\�\fM����qY�cGr�?�������@�W����:��7[�zȏ����{�N�ND�v�bKT�
{���=��s,�{B-#+�Vx�Z�%��/�(?��9&s4]���5���3\>�P(y
�6*���+����&�sN}wT�$�8���/Aa�ԥ5i[����x@�� �`��������4�nc��,��R���1��q��a��­��[C���	�~n���7a�F��G�S̻1[�#ݹ rŀ�}�uNʂj*�6I�VU˕��UP�����h�1G�2�Rs���Ծ�y[�J�梵3d������A���i(Β�����~\@?�,�8�(ݙ"�i��ݤ�܇^��g�ms*$��ESפ�#-
!���U	�����lQ�̵��K�1u)�ױ~Q ���16������	���8@qY�&C��.:!�6��;c0߷s� ��g��"HSK�P
��10ڂ�|���}��([��`�d>�*��I6�c)<���H[Y�ғ���,~ �lvЧ%	Y�m�[��>+�8U�t�@�e@��v�AB�a������m����p��_ \�**�>j۪��q�E'|���s��}��)��Һ���w,���n�b*� M���1?VPg�>V{���M�|j�:`�@�������x��Ox6���Q���s5��I�a��P��'��C��ݽ��(��/(���Y�<x�̶H|�d��kѺ>�Y�G`���*"�r��l��$-.���A@<��E��u�#�n�����,�=�bB�B��^ͧځ[�<C��^� ��|�C$S+��G���.Ԟ�*��� AP�	�oe���W�\t ��i����� �D=CZ7��<���?��1����m!�����;ZЮ��|�-����;����ٱ��rO"���_�yF�
�`��!�;��U��X���t��(�JW9�~�#&�M���j�n �I=�x)��s�Y��rvHYF|>zBf�؉P�":�m��'(����n�?0 �捻Dr��Ox@{٭�Qh�BU��_FQ��(p��
�zk6=U�E��+��2p����v�)��Y��4`�n}��Ƕ��.E�Tes��q�e� p3I�k	Y�պ��ľ̫�}�Q�@�i���u��<��mЭ�6�e@x~_�"^X��$Ԥ����txY��&��_�/薳�q�1:z�3#9�Sd��V������#�����m8./����V+}����� ��jm�*~Ԉ`*P�,��\aK ������=}�������1�c,��s��E��J��3�2doR0�e��&��}
�)@h��}�G,;�`�͉BJ�Q��ib�]M%�%ᖝ�$�3���0f����9��.����l�O�u+6��,w\μ���� j";+k�Q@��7�HDi;w��d�N�Ž�͊�BX���+z���I��Ӎ�R��2��q�:�r��Ť ꛕ�4�J�\Dt��>w&�����Q�)�,m�k�b��	�KM�PA9A����C�T}�v�٥M���dҊ-"�Ҧ�^���o"�.��Jf���Q�^#��B6��&���(t�f�4��g~yŪ�Y5����A�Epq�3���Ĕ'�Д��*�AT:Vb��|���-%�uw�e�I��UU<��2Pl�SF�׋���t���ޝCɶ]+�7���Ld=>e�_�T{�+�F^Tx'M����DE�o�-l���P�G>���Ѐ]
�?�8a\I��$��B�Aِ�"�n��P�j�����Oy��eDH��t�k#�AX_�&��O�-���T`g��JK�7J��"�Ÿ�(64U��]'�YP��D���я���rZ~�xy���uu$|�2���d~���a�sa�w/���������&���5#k��'+��}PkH,h�d��v���Tϴz��Z��G�_ZN�ad$	c���Tx�4�nʤ��6�P�����ʞ���|�uxP�[�+l��VF�߃)��k�~1s��Q��"���c&�,�Ƶ�ͦ�X���ϠoC��l�I�v�$Fc�I��2!cY����RI����-䋴X�Za+K�k��Z��\�=�Y����n4a��gT���SQM����܁G�"�]������ ��wl�q-��/\y�u��f�ň7'�
�l6:�9��#�!X�Ě��b�����F����w�:N[h�[�n���=��C1;����M9"〧����;/Quu������� ��N�ۖ^$b����|7���V�Â��a��s�.X[�H��M�K/�evTv>�U۟��gSǄ�E�|���Hr2���}U{9��y,{�hh����y� h9��&5�Pg��X�s2� �b��ͼ�tzer��;�4O�+NfpE/�ݔ��(BW��r���9����(�oB6������픴Lq�K���xRtJ�?K((2�~^>��npM��Y��#�)a��ݡ"�#�|�a�*�*�j���[e�G(>�D/��(�|y�W^ x�m#�]���h��0T[fLL�j�~Ԅ�jo�u��9���p���r~��So��}�'�ť5^LP�1��
IJ�p�C2�����IJWC&� ���/��\���=%ݰ�){�����{8�ގIR�v
�Hp*Mi֪�X;����SAe���x$��V+<�$���s��\~�z�}x_a{�x{���#2'ͳRl"�/=?�z`��V��s����8�>�ȷ��k��*98��е��zy�i��S�h�4�?_�\;���Yմ%�V%��b?�����ܕɪq�ꑝLO�t���RT�^d.��p�*�> '����'b�CU/$mް�Q�ql�[�3@��pu��ToV�@���Wz$�jIgg.��]bT��$%
�?�H��4(eh��Խd�,�m��cn��B��
�b�9�uLT3��	yX��a�*O��;۬&����Ⱥ�6Kо�S��`�\�˙o�
��Z�d���%�����隲��/�@,���z��҈��I��cW��f�HЈc���h�|���Z#��Rt�Kj��N�\%�����n{(�ډ<��3�r��AI��֞��C����Gz�.Zm���J\i/��I��)�k|�c����l3	]݄K����'�q#��+��?_v}c�1N(��ߡ��~5�(5�T�Ӥ�O�!��n���0{HMWǥ<�����e��ؘ298���i���|IT�VDb�*y�>w����$�Om�~W�z�n�W(���r�
�z��Kȯ���'�q?Z�X���U/7���3c�n���e�����հ���e��Ym����� DQ� &5��}z)t�ȩԻK����k<�q<�2�1���<79��������8��в��u�F�'Z{r��(ഏ�,5O�o�ܙ�v�ʨ���Sn)ړ	h:ͽRj����D��j<s���Y�H�5R��z=�B���㼌��a�}���UZ�6�@d5�b��	��sV��5�n��7n�:�m��!�'u�	l��1*�Pte�
(���l��U��<$u�{�<l��F@�O���Wyl�@�+,�)����a�
e��k���O�X3��J{n6�Z���G�6o\�]ʚ>��R�,�g.����{Y��ma
/0���U�υWcnI�*%\��W�+�V�`õ�x�����b"�r�=�\����Kmk�)3��g3���	Y{�D�}<�76+7Ŭ柕� o�|feQFW�C�:?��\lS������[7tُ`@?����چ���� }zY��E=	)?YQQ��-ח�q��syBk�S�3Q�0�w����`�ӷ��FI�e�c�B�g�Y���_���x��l� ������l�MҦd� v��q�P�>@_�����^ZiE>�)>���K=��*�ڍI�t/��.%S�B@�����T ��/��GJ�{�fm^ͥy8��ro�Vö�ϿNo����i���ѓ׹F4�6�>jY�::�zֈ�K8�Ϩ]U5�SX��k�<����)�Q_���ߙ�%���sY���}�Q��*��4f�d�Q��*VE�z�5�
xI##:@�t�}��+�{�;��$Mr�J�������/�\��1x��U1y(¦}]ĤwD~���C���ڣ�1��H{�g�d��4=�Qa���M��QZ���ը��fGR�}�\��8Ғ�q��}�4;l��/LoF#�T��7����֍1�ޣ���'-�xT�C��h*��-'�I��M�ڈ�s��/�_�{�����G��L��z�����,�+����F*�޳V�����>S���D�Rg����;�m�.V<�����3�t�`#����N������M1��nܩ�7��u&�]�{جʦXO�k�௛:Rg�L2�4�Z��O�TS���q֟[� ���]�h���uj����X|��Vmwa�O��D�����K6}���n�Z��Oe��b�u��2��A�:vq��L�J�� C"<��Z��������������;��X���H���[���jB?�ݧ�#��Lr
���-T:�+�D֗��@�E�ѣģ�|Qgp=��F�uK�ܫN���Q��� B���Ƽe{\[7ҵ��H���n5֎6�~�b�.bצ�!�P�	�	G���k�눸������J�|������^B�^�Y�n����5��f]$g�(M,���D�h�t`&ȍ�f�j�7���xYg]�22X_7�����=��f��7*qKn�ֱhUr�Y�}$U��G�e��_~�T�1�;��j&�>��!��I�.�*۬�=��(��0T�	�GU�Weh�7bTQ=5�8�n��މh�\�_����+D��YZ�wr��V1Mw^im�G��@S�ɚ��� �w\E���Y�wStH���n�
H����v�.�ѥ�n�]Ux��D^����ї��ox�%��!�����NKx�#��:LۧYf<�0�W�z�4	ռ\agM�*�L��2�^caJˊ�:������Z�&���DS�zu`;%4��P���f�e�`�c�wH}�*6@v;���9_�ġ%�]���gƷF���S�T��0��o����� =^=�
���"�����P8� �ױ+^���#�3*d��T`� A���F�>�o�{�҅W=���ʾ�3�yq�z\�S�Ѩt����):/���G�*����fZ�5q^�3���XRg��X?��p�O����7p*�̄\���-��d[�P	M(�vQ���nS8�Z���j� 4!�f���&N!���[>��^������c���
��Er����ֻ����۠����q�c�]G�1}WUv仓!TE��d�*u��㴧����ag�1�Qz���,���R��yI�u�(֫�^�6_kk���	h<�"��Dk�y���'�ߋ�n�)�k�K�ngX,�h�{�]5Q{�q%��:�Dв��^ndH�P�m�R��
�>lB�D"�tf�����^O3�e�z�stX�g%����u�	��<�W<��m�Y� CDhkX�� ���fß�| An�G
�H��`�h"���L,���;/sC����HL��/�2mnM�� ��G2y�d�of��;���>$�����m=SfM;��&��n;	�,ů�)�Nl�]��3잡�.[;;˦��Ť��Φ=w�^��i^���`�#I������X$���}���L���l��4
��~Ti0�l8 z�Qٚ�(�~�y��H�`i2�>a�S��U.+׸��L��TO��<��u�@����#	�m�s��ӆ�u��*���~��fj�6���>�H+��m�8�B�������l==F���t��'Y����eo���|��$��tT
n���W�k#e��ND�\nB��.�l�,���=K?����p�|[��5��O �x5�L��z�L��Z˹H������ׁ�3�F�Q�Mr���4�4���2k���m)��4e0�$KufN���'W������L��3��̡���i��t��nQ�eJ-�X*\p.22�	`^c�9ν�z,p���ş Ɉn�}# 9|z!D�!J��W+�g(̏���\w��>�����	�O1���.��p���׹��\�h�(6�3��d'�jMk�XC�ݺKc�E���$K8s�1����m0�# �
�Cln�#z��gI@�gAЅ�t���:�g0��Z�2���	�1�6/L��%���I�(.-�}�g�
�)ޔ��}��_���OrV�^���xK(��Fe���^��"6�w9=��1�k�k/s�bQ�1L1ԃ<�)�N������uac?�{kQ���>��
@������R��m+q��j0ߕԓ���	&�Л�軣����b[`�����\�:��s	��G
�� q��H����r4K�;@��]	�D�Ӹ��$�����?�	W.@���)������%Eg��G&�Z�ɫv!%�h~�=p���~xjX��(�߲^0k����W��/	��kмj��P�
ʑ��Sv	�E��1~��R�)+L�
Y�� �P��E������=���WH�zq��{�3:k#� 
<.���?O��H�v���܍�M"r�I�c(��A�5�Ŕ����،�z٣�B5��~��tI��t��X�}�|N7pf���M�ڷ<fțP^�̙\}&�"׏L�p5
x�R�1yQBxV���v�T�%+�������j�n�	��E����#�}�z�-��S��G�=qN���P��76��2y�ɚ�����pQ�XW���4 ȤhS2P��+ZK��s؝ڛ��o�'���g����l~�`�f8)���>��z�����V��������?O��4��o��A�ΐ��&�d������^$�0��ٍ�47.V����9��B��OKH��<*S�����Gy�VJ��Eu8������\����)���kYp�<�l������'��|ݻ�NA~�ֿidC�量s�Tiy�E��r��x�?>W�F����N6a^����}̶Kn��
��-�����>��ݑ�O���ܡ~��3� �(��p85C���pR�n�{D*�Y�`e���zb�1�L���a�Z&�AE|�/Q�%н��]�d'�� �Vx���X����9ݵ/��t���n}"���%c�^�����u#}tD����@OK�IT���͛S�&��#7E�bή��>����գ�$?�o.��Y����DYP1Ёt��#��d �	�F�7�o�vؙ�s�5DZ��[ �w/�E�j�A�y����xR˚���cGe�����rO�I��d���r`�#��7�<Ʀ*Rv-:vE�ُ���?[��N�l�`0��_�����/�����4`0�Rp��3T�z*[�'�L�:��{e�]���z�	��*���I����ފ�j7b��~�_	���8�)��PV�z����D��8����Wdg1|�z� �(�߂]uB�p�:�%��dS8���Q�B?WE9Tt��̀	�ǋ�v��7��,Ö���ip@���ڷ��U�s�}sk���c���;���r�>l ʾ�����K2����"\ف�{>�!3 E���o�.����7��D��vv;��Zu�b�&(��_��eD�>2�H�TA�E#��s�"FhAb@j��%Bm�@�Yz��X��'hN2>��������M]����>�T����.��ʂ�`���<!`B�ju��`5r���`"��$	˔����T�F@�m�\�(k|����;c�XS�D*�}{�!ODC!�x1W`G����a�DG�z��B0�;�]�!� �q�F����?�8K�I��0͠����0�C�0\{�>�'@\�Cȕ��P?z]�*�1���e��C>@2e_���(U$���#S<0N,�t��i�;������'z��'�]�cDm
D��#+R���_Պ�����a^�����J9�
S��%t�p�������9�{�F�N�ǂ��;=�?����_E����g�Z=��;��4�2 ��)��\~����"36�(��C� G�)��T�pN�s��*?O�͂�rd�Л�_&Ϣ�{���vX�v@�;Iϻ�^��tP�����p�?�CG������+�D���o�s~����~ߩ�Y0�4��  Kn	�T ~} T��a��u��J��}Wn���NRVՓ�v��#]��9ʂd]�,Z���̭L Ț ������E��,�/�DM�/}j��HI�O1��س��m����N+?v˶	o�LQ��6�W��@\e�p��uZ2+7�&�����~!OV3�\�Q�c�0۴9����wN]C=��%2�N�b�|��ׂx;����t�E��4L�+��j�d6�YO+n�YUMP���ɜdD�=`` TΙ$(I D�5��^8њR���d�e�ɰ�}v߸п`Q��?��{t�LF�/��k5�Y�#b������&� �iw
:S���\�Q�vQ�a�(��Ͻ.�%�X�z\]��J�K4��}��<�ư*9��isx����?{�㕙* �(��z�׸��Us��:^��]V3�M�߼?�g�皖���rS���jjS�s�g$�e_2'o�G$�����I�w^��'Ӻoh�"��^��W0��rK##��9;y����܅,I� E�ӴMa�sv�!��?�t��� jG�7ښvD��΅�����t����s¼�0�������f�t�7��(}8�"�>�����7��fTP�Y���ٲ����A�T�t�]۪�pq�఑$JF@�@m�M����]��P�7��}���˽S��@O�!�ҵ��n�׹̈́K��X&)G�m?a�S�U#ah%��	��(��+������Gyw4�L7�E�;�r�\1W�}������Rԉ؋����R͚C}Ύ<���:<�����q�\����	�d
+I�~y�<xxQc�F�&	1j�6J¾�8���,r�z�]�U\Уv��.<�M�]���6�����I��B0�a,�[-�����C�o�0�qcè�����t���m��y��`r����l;[��j�7����_�:�����°ԝh��l�k�^;�� c�eIv��9�~}x=a�{R!w&��ݒ��b��v��gO�����\��:ټ�?�[Zڱ�i�	$H����;�\3G�s�k��"h��]3�oz�&@�NV�	B(����s8�WuM���؀zw��(eJ?����,͎ø�o�����1/�ʙNك���A�]>?��bby�H�������OYjŝ�.~M($k*���AD����9.Mn�w��sۭ;��WJ�u3�j�o���� �8]�Z��Ͳ�`�:��� �1H~kȃ���h�g~ã �m{�xJ�}���f�;_^ܽ��<k��>m�&p�h�������1SEi.Jƚ� |N��0� �#�i���_e����{+/"4jS��O;>��g����rAlP������/>àÛ�Rʓ�`��r=����*�U���G4��_fx�"�Ǳ\�X�A�9۱n�5���1��kЎ��y�-��9�1t��&�=�����hN;�}�.~7o�qU�+��照E&�V8W;Ͻ>{PB��ދ�z&'�������	���t���LgO
�,�9?{����@��`�7��������!���[�ʔ��H-20f#!)�99R�4]���IQ�T��f?� �o�3��>�%X0{�}�R�2�GK�W�5�l`o�AK�4H/����dwh�>-�)��o�C��.�r�C�f�����^�b��,9Gc{,^�9���9�u3����o���&�����j������-�T����،�=���t��������`�T����=q�����bff^���@�ԧ�m������_�ܱĂ���H���vr������=�q	7�Rg����_I�/-����|؛�>uɯ��BQ�o����Eþ�e�����A�!�;<�uz*}�wa�N�����&wr��?ȟи^�v��`��ԺP��͂�OB.�,r���	�߲���q��9�?;�Hs1��s��#�U�Ӌ��*��2�o
�n綱� �7g��J�-��u@M�q����"��ׄ�v����Ղ���vW�T�$������S���N�:~k�m��Tr��X?M��nU����a(��̅��o��i@��[����pj�rNpX��W��?�h�2�2-���`�W��/��*����؜Ps
�8 �� @��ݙ_�c���5�FL����;qA>� �k<~�Y屼�G���ōv�Y�7\/䃧�F�J�8O��.�Ҭ�w�;^���ӥ���64_�����
�Ƨ�g�l�N�]9�z�N$Pn�v6 ��ƤK�@���PZ�N����fM�*!��}]��`v����

 �)!���2CJ�����L���Ӭ�>��뭠7���;����@��egXa�3��ay4�w��)��/|)u�4��3��]`c4��<Iٰ|ԩ��T��Z�#�l���q���^�������<r�3{���;"��
Mw�����k���L�j{���i1ڕC�ch�3J6[�#Y�
�o�i�f�u�Z-�@���|�.�g2��L>�	����ʰX������HreA_�pw��[&�����_�{�Wq��pL{��U�w"��RMk����2�zœN<��>�4,M�z�B���~"�_�z|
j�l�T��Q����?{4�����~N�_�ƢE�v��H���ϩ�#��GO��M�/�֑�k�.H�s�>\s5��I�&ڇX�̒��g�0���u]^;��d:�����S�K@�#L�{�od�F�,H���c�\1sZ)5���u}�{B����L�5�?�T#^�:G�-z�u=�ь�FG�C����s�u��j샱�'��|��{���C���|���<$11��];����#Ъ��]4;�V}s|�f#���|НS��� ��m�J(���t55��E��8���K�=�)N&�}���U(�ׯ���w��(����;�%�RWu��J�Ś�I��~��KA��;OV�@�~>���TI9�cz ��*@���򈌴(��	������{��Ps%�n�E��轶g�;*$P��U9��5���_����wU������޲��*�w߬�P�D"��f��"��\v���i��T�ſ�D����'л�?�?�c����������!��*�r��Z۶�+����8�W��N4K����0��P�=A�Id$u�ߪ�-�S�y���m[�aT�����Kw��x_�ȷ��j�������hg����=���������7�0�4�1����@48�Iix��<$���1I��gb`/�V��R�l%��'�H%F���m��=����[��=N�\|��(��	/K���J��γkpۆ��ew���&��r�1�Z2���@`������lbj��/v>��y\m�@�J�0�,!�r*o��)<���QqaaÝ@	r_˦K�d���$�����k��m�=7�8�a��.ľ��S/�F+d�d��]���_���9K�9�ڼ�KO��D��sh�����=}|e[�K9{U��햲>���v���8�O�ʥl�U[�Hx���$��Y�/\��Y�$N����F�	}}P�!���==2�:h~]����y��cQU�ք+�5����LE礮ŭ���
�&3���O�R��u���`HUE����;��:(2S0���1�|�Z�RTW�[8{0M*���+Aj?���!nm�4��&��9���CO�ZF�v���|��.�^�kz=����V�ϰi��=�։R7�|�!hR�� �Ra,�7��&՞Q˺��.��#�vg}����2��B"4C��/�̵4�}�QֻXل��%oj�@�������h'$ЪX:p�¸�wh��	���t�'/e.83}���<.�;���8�U�z�������"���==���ӳ�?Β�:+���=u���oS/������U-���?ǳ{�)9����:}VL5�)���^��.��Y2ri�g1~��em/�{�ȅ }ȉ\�����ޤ����� ]g[�M��޹ժ��q��$�)]����(������)���0��j֧�Q~֟Y����A�yוGEwThe1/�67z�ظ�H�J(�''H��t~Ş*���Ҹ�ϰL�̐���!U��"�Y��f���g -����2���j̞�(�p��0��]���v�z؏X\���̫�=.�jk?��[W�V��o��C})M2_x٘��-����|1�<��JU��''�y����h�P�W�#��������bvM��e�����ְ��2~��N� ��M��F��ͩt����ʼ���F���U��y�\Xp	�Q��uչ�0Z�*�nԔ��;�!�k_��CN��x�E����PM���<��i�AՓ�"
����E����������^��7-�e��ƙd9ʇ*��x��JcJs�>�ԕ��M=�EC?x�#\I�g��3U�{7&��f=�Vwh� �l\l�h��t��+��
8��l�e��h&���7�<���)�'�Kf	����ːDz�r-m�C*d�dl�ou���"(�bV��_���d�#��a�4�`��O��%�lӑ�:
)����X�B*���������RN��
��sƁ��� x�)�+�����.G;�G���q�_����F�(���G�~��>�~_&�6��0`��(�[�\�N݂]\����t�?����s7^���//��s2�PK3��� ����C�FC���K+]�)��GCi�H��tG
���&O�ݕ�bֽ�:^��6�R����$�Ԇ�Ig�g���Q�ˣ�j�W�OX��W<�����DX|�����Uu���qu�	k�Je�Xpӕ9��)�d8
�Q�a�9"=g&���A4��wL�|���g!W�<�fJ����oh@|��|��N�`w�;{�>�r-W��nN�	�M"�}i67���#Uvß���+����eI�~�]�3}�eC �ؤ�qc5�
Z�:�z@��5(.�Ƥ}k�Zs����J�?1�7k����<�����xf�	����^���$U��.�Ս�7���7��q�gV�g����t��Mgߛz���j����Q�?:��������;l���0�l)�J@�@X��'��jwx��پ1`��p����~|�<�	>R-��鞬G�M$�_x�i휱g�i�
�7$ cE��ɸ~�O�T�L�I���o_����´�nI�y�/$J�L��ȆA����2�׿�F�GF�=�I	��a�_r˟ ��P��j��3��q�iL�N�����$��/r�J�o|���~��bMuuC��E���%�[�*R�{�����ĭ����c���όI����K ����u:�45��i㫴x���CM����8V/�,1 F(sa����j}W�I�{ZH@ڃ�NL��zxA'9��p���PJ���`|ĩ�֒�h���CO����t
ujL��Y�7�a����6�����w�o�x�3R��J;���t��h E׸���z���7�KX'�x��ڢ�ULW������ipw���x�M����^]��;:E1�b3�6��t�'�OB[�0B_�i�6���,���Y.L��y�ܙ�F�ouZw��O,3$m�r�}��6�>Cx#��t��8�����QM/_ߨ�c��X�
�DzWi
�;��^#��HWz�{�� ��.%AZ(!�����9�G|����u׻�k=�יٳg�ޟ�e&|gB�/�!�>��	[�^l�I��۔��<$� ��rŒǅx
-V�-��T����T��h9�	��oXi�&��I"���yEH�;~�.k��b��MԊ.l��d���u]���m
��3�����8'	�Z�s^eh�����<9�hW�!j�S�w+GǪm����o���%��#*��x�������i�]Sr�ytfh<Y]�4��i?O�R�/h�7�$]��ث�f��\W�=?.-3Z�X��e�.5���'��8�o���7�zj�3_��g�E-S�a:k;�o�3]�Q�j�����������&�y�b�kJ�:%�h�R>��9�!j�+���� r�)��(�8}�S�۸np	�}-�hI� RT�L� ���<���fH��n����``դ�+�r��E1l<��
B���LrB����G��X�c�[Hd��<6�� �/o�M�R7.u�����qt�i��ǰs�3��\��h�#��ʇ�]�k��|~;�L��y`�0'�D#�L��J�""*��#r��6)�^!k
�����`O�Y�0�m�[����Z	>'�g���])7)I��\��6��*��8jO�SjB�6�ȨUW�m���Z�=��6-g��X4OK��K!i��@mx��=��:@����"r��CE��"��i23n��FƬH�S�U�Ca���m���Nc9R�i��,2�Rk�4>�y&���H��^�OR��cl;���*Z
��Y���\��&7�X�s�@��w���Yw�~ W�Wǵ:���E�B2�s������m��#��jz�}���rV)�|+I�յ�y� ���7&06�5}O�U��/�a�+�~�b�m_ �f'(��޵_i�OR\n�@`K��p����>�ACf�d�<�j�wgC�_���B�)��6�ͯ�ne N��_�FA�sRG�{ô��� >Qį����U��:s�zOp����551y����8́�����G�������.�k�5o&���(�Ɖ&dd���F+�q�=�Y�"L_�G"2,�T�嚡�'��ܵ���)p�`��p*o�C�EB|s>>���!}t�挿����qZ �\���mK�W�G)��|s�Ɨ����s��k��s_���d��#�B7�1�
lBR�EH�u
�|���ǝ�Qe���%�Ñ�u���J��%͸�4��O������~�"�͢����#0�OHK�ǃā�8�ǀ^�B!}S��F����Ȭ݈��j�ykG{�A�P㞣x
�o�USu�Q�[��ټ��!�
e�T7f�<bM�īvk��ZȦ׀�Ɇ�j�$2��N��&��ϛTCۻ��o�&�k/���u6���[,���6!�2BjK���x@�轅+�,;�2ʻ�n���úL��ب���:O�Yq���5��+]}�0�b>M�[��V5*VRɄ/���ARՈ��o	��<�v:|���`ϰ^Z�ƹ�I�C���ܝ�:�TY�$t�Qr)��}�jM��CTS�k���v�1�諸�[�b��nv�;VQ�resK]�\n�dG����'p�b�V�L����k��m��_���[n]4Wh�gGi8�"RW�h�n�ʷ�!���Ş�$�3�n�w�-��"'��4��o�	�YWB�H��#�3h�D��_�mA.���9̳%��q�Cb���{����Xrz<B��f!��E��[+tX�z�(P�rZ�`��z��*68���E�m�NY&����n��<a}�(�j��Od]KA�vN�>�e���+]�
s���'*vP+�>	�-�6
�[d[��Yj��oh�*�кT�:z;�38߲� ���ƒ�8k�vW�7g��[�7B%�c-���M�M,�*�q�L��.$��$�w�?���=a�Q���5)�$�
ۋҰڞ�}��s���lU���^Dg)Ќt�q���[��������)�&�>��K���6��FrY�`{|QU����=�20
 �*6>��$�O0=�U�Mbّ��L1%ios�<p��l���ot6�m���oI��V3b�xҠ���W��Ob����A未c�[��zq��8$�����:Ӭ��\�o��Bܠ�z'|���I��zẶ��[��5D�k��+��
�J�'W4�����yߚjYE�l�%6΂��{#��+�_#�{�?�9���X ��}�U���n>g��͕�x��C���Z�~�9��ۮ������DX;h7��wH���~�@@��d:t���@��%�P���i�Z�HLLY<su����u	�⮦1���}qa<o�x�9�e�?n_�|�RQ�
�gT�>�g9z����j)@m�T�V�]�l/&�~�r.�*�A�{#w�dլ|�:D��+��T\}!��³���#j��� `��:�$k�ڎ��>0$�<@s�[�9}q
�K5M��$�y���"�'�k�Z���E��M��|c��:��+w�e�@�a|�;l���V擖�:]X�b>TVw/�2{��)��5ta��U����.�k�3��w<���ٓ�ҜD�1$��σVk���k����-�{������#h��6�ŝ��LqVuSU�`kN{�嚰_�M�.��}�@}��ul���Li�S��g���5]�+�-��`YTu��x2.��e�̐hY2�~�=�j(���UU-�7�&|����Z�"[�%���dt��W%Me$��ɒg>|��U}Q���h��{�=�4G_��x%�1�w�^��R�Wy�[�̩h�h��B�[�B�U�r���Dҝ͞��V��-0"(vߍ��X|�����*���*�l�DS���d��Ed�L�[�~G;�f�Z-�ж�%�Ȁ�|�>�~�@��Lh彈��6z��Ͻ&	e��J� LOot�:x��Zg�Ϟ#��(#���.�Y�L[� kC�ի�.������|�륟���a5m^�:V��Q�T�c. ���X�	�BϹȂ�fe����99
/���YZ�h�c���Щ��A�ac�fӢ���ojA�_�b͏��������ߞ_ ��z��I���:/ r}�,��C "l!w,d�{q|��Ǟ�������sVα�m>�Z�D[�N�85�
�m<Q����)w�������C^EnQ�S�w2��X�D+��J��0�Ub� ���Ė�S��r!-f�X:m|×/��R9���7ƽ�4u���]�&�/i���Ѵ�>�`�rX��,�,����q�ߏ�����jk�4�������$S�t�Œ�����o@$�q-��L�`6�L��Aig���gc�ᶂ��p9f���:�����F�i��}|�.��E��+�ɴ��[}�!�377!V�W��v� ����(���fūj1��i!S��w�x�=x<)���!5����~U���)Db�[f�:S�i�4�+Ͱep[5MS-[f;�/-�4�S�mX�g���e�8��E�nIV�߶��<�IR�D�+��s�
H��ZU0���Q�㙹��%*�D�r����-���G���w�����׊h����a��-R�U ^z/�_-�]y�e�8;�M���+_S7B�4�
���Ro�y�m�+?	����\�ݫD*�_��&���NI)�;t��&yñ][+�"թ�!y��˙�z�Ֆ$YC���0�e��[|ح1ʽ�y��OM�zܭ��|q����VΦ{U�Ѻ�z��֘��XS��y�"|��;�i�x c&3�ڷ��k �Oi��[ׯ�6�m3=?�U4�ݴu��x��#1�x()=ׅ7��'��B� ���Y��idr`�X�oH����5�2��=K�hla�h�l��MY�^��$�N������Y����*�� �R+����-;��ؕ����kƱ��[9���{o�XV(����P0O~����NV c����r��S�E��"�6���@����w��Z݁�#"]�b���)�(RazG-�UC��gp]�9%�dw�r^)6tt��pҷ� �7��uX��g)k�5��q�x��G�
���6����^K���x��0�c�sQ�&�H����a'�7{R;���l?��X/����
Q�^*ik�����8a^s<e�" ��N��-�9�t��u��!P-�����'�CAէ�W&�r�+��f��]�߇%&a�k>���>֯�����JW���U��Io�� ��^�������޺�ni�o��t�_T�u7-����C�$�H�l�7w`�k����Q0 S�[�f��~��I�\��Q��'�6���L[͕6eE���*�#��	Q���3�R?ې�Q��"4[�3����ʘ�Z���eM"��\����.�4�\E��s;Q�i~�%X��X��@�G��?�9e#�~ �N�DV����X��&;a���L�)��6� b���w�9�����:��>z��w��7���C�5�&_@�	iI۪�|���F=��lG�2R޾�wyJˑ�{{�̱O�_U�S$z�3�O�qЫ���{���E*#1�x���P$G����GƄ� 5�M�'�<��|����9�SLf)�Dn.@K�׬�D7o�Љ_��6`6�^w Չ�� �2�+� �D4��(�^�m������@�᯼E�'��C�șq��d�Ze����D��]�.�+����:�t��ʐ�5�>�M�w;+'v�pX�<9O�������r-nst�o�Ho�P�����ֿ�<�H�LW��Z�eN2��4���O����ؕ?�{?�id���;�9t5|�0��M����'!�O~���ᰣ�	����E�>����)c
KV�z=��v�cv4Qm�]�%l{_�/���J�z�DԲ%�������T:�G�� ǂ��-�k�=p
�h*_.cr)���b���n��B�����M����ŝ�@7wT�
�*�u}��ļ�>�Hnd�m-��t�S˔`��mX���?'[ǭA�64�3Q�E��u8Έ~t5xխk-h�3��	���f>�9�r��i���t�m�W��x(��;N��&���C�ig�L�K�yeMHJ�7+<��T�I�������U���o�,���[U���@l{�zh_+��~��y\T{�Z|
AA��S$:w��	!�YUa�|�u��C�^U�Ms�����Z�Pqc9c��V�/�a)�
�~�F<|'�6%�jk�)��@��v��x����6�E��EK��+�rx��u|PH�	Qq򉶵�{�T����O�ԽOڵ\pL�Ś�%��S}��pKqE����'	U��8VP�s0��\:�T��5�(<��'�K�Ι���5.�������"��U\��H��"N>X2��f�p
[�e9� OF��4�(ܴ��ͼ���)��t2a���(��R]��*�
�2y B�0�,�
�I/�{_/��bsw�y���??~�U[a%�3`+��կ�DU��ǧ����>��1Q\��
�l�����<#u桅'�G��3�������@��:�[��Q���a��N��м}�Ĺ�*���&W,���.�8Җ|�t����%U�Bk;ij��gpM�̅�v!)�\o�g*���bm#I����a������P�!;�X��Qvn3OU�L<;���tENe�[�@fv�p �%��s=yd��ѥ�~��]�]ҹ��N��k<YZ��Tl��c1���1e���\@YL�Pop�R �[� *�솆C�XS"��R�O'� +?/��$���U����N�z詡����-�Ƀ�-������y�z ��`o w�ne����~s�>���2��Д����R��+K�M��]��tų�Ӽ�%(ķ,a���5)n>5ޣˡM���	>��4���;��N���R���2��R��&�b`�\� r,s�����e�$��D2�ɑ���jUG���{i���XOmu��[���T܋�3V��%_ҝJ^�:K�2�����ƻٳ�P;\�~ϔG�)�Н �|���R�����m��r��[W꼟�Fi���ɯ�6�|�^�^ee�Ʈ�trL~'�݀���ee؉)e%�X�����u{}N��:�!��l�4��n�c���b�܉m�?��CN֖̂Qq�?��@�^>�f�&�ȃ�[o��M�B��M�"xj�O���l�=�������ǣո��x
�iǩ8��|��s���׶8iw��L|_u\�����c�"��il�1�>?�*5O6O�@�����H%r��M|P�6n;o���-8�BK%_	I=~܋�ۂ@HSVAeU�LV�򛊷�y��t���=ҫ� ;_p^y�T)|Y-ϻ����\4!>��z�B.�|��҅�<3{z��Psv��Y[�Ϗ� �L�6b'b��:ې�싮�,����=���7�$��,'�1w$ׅ����C��6
@�9�J���F%Bt]u�*�+���4�#@��߿t��*0�iZ��!a��I�VjOc�т�qq�K|9��'�Q.4Wڐp�~���D��9�I�)�y��N�
Iic��  �A!��n I�p�`�p��[q��9���6�HV��`�WF|	AVMw��/��H� �QTJ@�˶+�Zt��5�f׾�y����8	;`��H|���a�zk����'ʧ처�S�v �Z?fIﭠ�1��k� �X!��e����^c(D����ߊ�y�E�A������F���)%*J�H~DR����K�I�,ѢU��A��;a���j�]��-� �0��6�%���YEb=xk��5�Bt�h�$��R C9���N�����ҧ���&Egc�)��7�:�(uaU/(=�H)<�ꂊl�\^����L�D��JS�G*!��Թ����6�U��O63T�����R�W��NIt�z�sڱk�`0�-3	 N�1y�S����3�"�꽡Bg�B><4�d{�$	+b�Xez���zԞ$@�	K��2���9�:\d^_�݃"�u,Օ��n�UV��Rd9��s`6w9[�� g�?l���R��c� �h���cB�b�������^��*�q��9N���*vLZ�������e"	�أ��Kޱ��$Ia*g%��.��9���mXj���/�1�j��@p��d�f񑈂�dʗ�X�S:�l�.f�w�e�u2�߾�dr�}�<(��1���k�}��sJ�Xm�̩J�.��`�GGr�ԉ��@����]3��������^LG�e��O�2G�n�"�� �7��aʬ�ry��7�ۼ��}b!�����Ĕ��e7�WW�Uq{�H9)�ޤ����O�b�G�x�T-�gK�'Bh%j�2��>i�����ȴ�cJ�/De0[3���c���p��'����ȳ�N��&���%H�o���3s�u4)9}|�=�*�,qV����߲{�+�[���_�L��XGY����d�m�nz�ƽ��%U��2�Yʹ���c%$��Y"������C�=�`���Hy��*�C���@���s*R��CDÉ���Д4��� ��9|�)��׿'I�.���/�g�}1���������,����j������ ������~������I����w^b�����^����?#���S�Bw`�������86�L�C���0����^���%���|q���9=d�4�+�ލ�l��!��]�dϮ�Y��5�:���-����%@@f[�J��'����@`�Z4o�k8gԋO��>�F��$_Uy��D����L���o�soߤ)Qˍ�1k�T*���Qd~����'��<����c&%>�:�=*�k�-�2[V�z�>�f^���4}'Xh%�3���Ĺg�X��~�~0J��d���po޶�ŉF&)�CZ�&�'H��JP}�<��f�*'ihV�����w���D�2����}����C�AA���Z��U���{�3��߭2f_�N����7P#:\�`�[�Z�ïa�8�}�+� ڟ�*��Y?���pMv_)��2�Gz5Ri6��t���:v1^�^D��lk��Z��$Iվ�WJ�܌�v^K��%li����~\�x㓈�v���(�!�8���w;�E�&�T�������
����Z�+���^��s�c�z�A�Zk���[UM{�����{�a~U}	�g�0|���RH��^��� A�|$�x�*�Aά�����"vW�n}#��r$Q����@v�&�4�[{���Y�غL����M`���Q$�|xq�xR���#l��#J6nf���̪�J����7�V��g{"���@��}�-|*�&	��|�y��
8����s6�����e2%��
����X��C��}�U{�T��
khO��
1���C����9�p��
^����:ع4O(�mJ�A��g���!���{���+�M3��fP�w�&�OG?�|E{Y(B5\m�l[��'��l����Zo�ը��
�����aJâ��K�M&5�-,��H���md���<�j||>"�>_�T�r����~Iq����[�}��Hy�(TM&�`��i��rGn�t����,/2R��!c�V���{��{��۲N�ǈ�@6p��&���z�F߷ �=���!i������S�c�2!��C�%Ȃ��;z�b��c@6X�=�j�ve8����4i�2sF�೩����(��"C�À����a���`�����pn�NV�H�p��C�FDD�33Ծ���h��AO��+��e�&���ѓ�)��|ȉ�B�rOxC?��D�����9@��햎ײ6��c'��y(9�a�v�hV�黎�X4d�j�;�����+�v�T�����8�#Q��d<���õ���-��C��&���cD\D��O2�����+�`��J�VP@�́��Z��!��6�juu���>-GkX.&ᙑ��0�hw�¼TRp��W �W���u{
,>MaB$i�R;2rr�Za岦HUϖ� 6r���-Y�tH�;+�e!�������wH�@��P��|V#kV�ݬrO&1���8�ٺ�Iص��$���?���o�lg�I��D>d"���L����hM�b�(˚{
���ha�\Z4\{�*4�@n����k��i�o.���8	[�t<��q�(C�6"��T[$��$�d�~6<��RL�(��Ob��)��\ �J�]CB9��e���n��,��4Rqp�b����gٿ���T�=C���i��{�l	�Qv?��Ņ�W��r_�C5��;�K��V4���0�ј�[�﷏�=�[�٪�����ǻ�Ʋ�~=y�]�9-]ћ��f��f�i�̺!�	�b�E�����(w햾�w�Oy�_iٵjﾹ;)���}|��8jt�Qvɦ-� �����OD�����gt�m���'�䞻����!'ݭ��ok���W��Z�N��}k�L|k6' ϻ��~�����銿P?v<j�J����?k��vtH���J��x��*D���E��.r_+^�����D���+���$��[f�;SvW����J����t���5�����U.j�	' �nw"6�@�����0�W���,�+>
2��씎E������	���QI���0��>�ik�N,��U#���p��r�p�ũ�V�}����o�������� 'q����,����6�kLW'rx��e�>'Q�u��j�����S֛��������a �7��
�t�Y#>��#�5}Oj!غ����ݨ*�*%8�U@Yp�έ�njg�ԝW���a�q1QG{/�-0'D��������/�������L�/�V7=^�{:��R����v�cJ�h|���\G�,���SSo��*��Y���d}���iX����wT��&�0��M����� ��U���jq�6eA�����|�H���B����� ������!<.���@\�j-$��%�^�9�M᫴/T ���ơ��;�}Z�Eҋ�V�9Mm��և��ߤ������TdDT����i�0��9�(�U���YH\p�f�ïL�<��,�����NU�1�bg�>�!�7�W��8~[��!҅���<o����}O��А�]�������i'����:=2��m�^�=�E���4;��z=W����t}���B��#��%Mb+��k|ޡ���	��@�PuZ�l�ע+Wv�y\�eWf0���:u�i��b*p�}={|2$ry�2_�ʊ��7���5��1��&�ۯ�����uK;���|5�=y��4�5x�B��]T��y�(B~TOA8��6���$N�p�ˬj@ZyvHh��jrM(b���i�>����(���-kr�TŖ�����u��Ğ��*��z}��k�6� ]	K�~Ř��p������=�.O(��~�[��Z�����\Ӣ/́��/�ii��yը����O��%�[A?�H�>��䞿N�%�8&�IW��ү~m�Sǁ/���ܤz��qG�Y�,Y�n��ք�zD�!�����e>+P��vʫ�~�=������T_�e�>��|�wJ�"��z`�T�+�;Ojգk<ޱ&�]o�Ђ싮&Z�2Y����D���)j6��p,*��֏�|(�@���E�?��M_�[ �*\����缋��zE
N6���s)1��6J�6�������rDG,���x��Y�Jջ��iЂ��B�|n�E����2��4,�iN�Ep�݌ii���T1҅T`���]���W *����oUS����ʆ`��<X����3 Xx�b�@�!�7�\����!�!�4��3T��hF�Չ�bx��M�}���i�K��+��
���<i⦛I6NCwz��m�v�F#�R�r��5����y}ҥ���7��N`�*��½���s�O���3Z{7+-��8��ֆ�V��Y��7<�i^��;�4eP�a�hi2�2���ᕧ���~J���<O��%�Q����%M`�ƣ'��9c��)�.Þ��Z�*NÞӒ���g�6D��z殍�:;b3�ӊ������n�e�秫����\N�`�9��������<v7���Ƈ�$~o�y���ޢ�:�0g�y�%0�w�Ea��9�^伛��a,�M���;���P�T�)�3l�%���q�>�S�߽ݱ�������]��'�?�)�g26�7���`���D<+.��ۏ�?��L����)���DN3�����79��<�ʜ��%�pjʤuֵ����	=�n}����M�S>�O5'���k�1v�[Ke�vkS�.�����ݺ�)(,l�1�����h�5',q\�MgX!U@�Ĭ���5(��{m���W����9uSS�A��������k�r	X���A>�<+�U@��tБ��=���̵Y�WB[͛�$<K����EL?ui]̺Ӝr-f����w|��*��>W'V5?>%��c�F����LR�u��4ۍTa;Af���G���*��n:�R¹/�|���8������[`u��$�-���,�������ӞZ�0_���� �RH����sԲ<�<���GaR@��y��+	�Wn�?�ʜ����%h�!��(�l.O~��Z��=�*�DI�]:�S�G�`���Nd��������kVb�&gm� ����'Y=�hO{Ƽ��}���N�X���
�����[�\�����?t}�V�M�0C���o�\'�>�P�?��d�Qʨ����1�y�[�)G���j�n��8jf���z&�Q�ityr#�Ϯ;@��IׇV���\�|ˉ
�|!�$"BWɱ.׆(Y�Y;+/�x������^���z2�U9�V;��m͸ں���Z��+�Y��8��>��-T\^��T��Џ�䝒cq��R��m�\�/�5a[]��m,lEJ��Y�Э�4�9�ǲ���c(����_Y��[�d����B�}v{�x�f��?���Q�������r��FW����䙩��r��`8�礭��kK
=��t'x���-�p���Q'</�+))Io��N���O�b��A/]����j'l>�^s����Jٔ�hy�ONӽ�g����ya�f��A�C����'<�.�� �Eq茈���O�/ӎ���%i���63�����e�c�~}o�>ͩ__���i&F<���W��i�;��ӽ��J�u}�6��Ox�衉L�n}���>Gu��(g�ޝ��[�O�D73�jڇ�����?��L9l`N�~���@�J���Ldtt�#�^)��� ���`ϵ��G����՘A�{~�]i����z{��3ix�U<1ES#{Ү��Օz�E�i$G�׉j��5��ΏlG��� ���QZ���B�]�Q}�~��Դ]4bc��X�s�����JK)X�y�ݑ4ϬfEۈh���Z� k�iJ0��6+J�~��I9�3�1����)������E��(�ds!F���pv�쌘5���^���y˹��4V@��f�b��#\�~mmm�di.��$E��/��;i~dH�'���kЍ�&��K`0��Ȅ��$v`T9������iJ�w���]nz��?�9�iv}�c_D#�#��� �:�����N�>���L��c8���Xdd�ܑe>�<k���MrV������P�;�݇�9z��`�Vs�P*�ƳcQ��=;;޾�5�y�.�;9bؔs�ڵkĦ)^>>#E£iJ���-����BQ)�T��Shcy����]�X�&L8��M����P�@�k�#��������QUMmֳ�d컿�q�<1������5S_jSߍ�_���@��5���1��!�6+�MS^�!�V����f�L$f�/uf��)�n�a��]�_`5ݹ��3�4P���:&s��۞$�#�7;e��t�5��\���gmy5�5k��$Tf"�C�'ݺ/�w�^\�|j����K��5-�*R�@�7ä#n,J�����p�NJ��� (l �!�TU	w�^7�t�KH`��l�%9��_?;#�+ ?6��N��g�Nv����u4����e�d ����uj#t�jCG�l
]hQ�A��陘�\io>0�244�Ƹ�O����t��ׇ�\�Ħ53X���1���dB��8c�O3��,�ç M���K�����0B@�!��R�GA��۪|Ǧ�� ��T��$�۲�w�G&� @Q�m�!D��N�.�y�Λv:���`0M۵��ݑ������@+��6�e�7f�SRRz�R�(�Gp���L䔖���!��e���?��F������FH<�i�|�y��n�%�,/�.�y��1C�-kdj�/x�HR�ABH+q2�;��}]A�f��<�:_���jW�/s 	hӯ�B߾���<ӛ,�ׇ?و>�ݞ@�_E�n���^�1����E4탊t
�O9�`�m�h4xm0n��]q�{�`聑��z穆`��mf8X��w����!t�;ݦk�w5�1?7�K��������"�[�SJuL���#�c4f��C���0W@� u��y�ޞ��Q~%�X9�!�~��+°�gv�k8T��y��<�"�i��xe��z����i~��>)""bfq�������ג$���`������?��������Z�ciP�a�-jj��s����Hg�b�e�8��4�d�FW��ו��Wk
��.N֗���</�{7���B��<�#[��wt���r�4�Hp�~oy��Yb��)\s Ja����a�!��K'�!�F!��ԿkN5��5��f9�~���fW�A�B����;�q��4��#���5�%��y�ɺ���ݼۍ������,.l��m����Gwc.ǜ�>J|� ����̧O�0U=����NN �0ź��Ͱ�wu��n��������i�����\j�+�9?���ܻ��.o�P�>|k��33\�~��S#kQ#���ܝ����@��XǫS��aL�!��g�ai��U4B�	��e�c>l�1|I�N�X����7�1}!�ߩ��s�{�������xえ��ʭ@w��&��-H�w����[I���΁?����.��~���j~9�k�_�\/�:�Fs Q�#{l���3���.����us��=dJ���J��á��GVN�WjD����"��O�?ן
=�ރ�0�a(P
Ŭ�f4�72u��F��4�,s6oJ�(�j�� G\�%աV$5�cI�'�;�� �#��A��i1�[_Hc��G�N�`6�N�W�68���!�� [�q[��Ą[� U0���s�Y﮻3��̑�3^ 7X8�:|bpp0P��� `�����fA̛f��/.��{_G�����:��*ۀRpv������	O/��A"1t�]��JO�ز]��׵�k#�#]�ă��*�@f��� �6�0��U�u�FĕK���~7����y��0`��r�գ�-��uu�&N���l�T���B����>bȄ;����*�s7���s�K-�#�K}H���V3E�B�w�q2�1��o�\��^�4:qFu�R�̐V��iAd2���%�.|p���S��[�}����AT��Lp�]�#!��5*��pM��Xp����#�rt�$���Z5~��>�	w�e���C�B>�(y�i���|�ږ�C��ߵ?y��[�D�`�(5�"��i;ފ��̯�@j6��i��V
��_鵌�Z�o�d�{W�<~���E�#h�l��$�\jTS�8ɥ���Lpв/����s�QGBنPQ�EA��7!�����k�ZD�+B-�f�c`޸��t�"o�T����'T#8>�F�
����W8S�����([U�F 8J������k<�o'�n`�����3��kߍV4B�Y鎬��ݻ�o��A��7��N�T-�F6���g��PB.;�*��J9�+r�/��yF����X��8���zn�T���G<�QA�a���ܩ�a��^��,��
v��/��sFiՇH���s��>�q�'+l�J|�1�d������B�xvv�DyVPa�R�e�0���6m���M]<uȱ4J�c���X���ɽ�eUs�dnGAv����p�� �R����9E��z����fEw�W�@��.�1� !6I��b!�HH�R����5.h��K�0;���1�wO�"À0����N�s&�1��5�F]�Y��Ai,�Xƨ���2�ʉZd�&F;{^���}iuv�{s�3Fri�?r0rf��$H[�0ȌX�D+O�;�B{��#�6[3�x����V:�@�Vz� ��:��X0�r��2��'��
˄*{Њf�x��	O�gb�N���O�t���7^~f��B�|���l��o����D�*�R����l��/�gEWk$��r� t�OL��˭�9����i�w\jN�\ҫPS�4�*��6y�`��CM?ɛi,B%$� ��j���oȥf�@���x3���#�;�Ԝ0�A-�.A'#f�VWW�b+���m& pU)�rt���f�I5�yp�<@r����� P�O[m�un�D��v����$�Ù����v�����*�I���f- H��v�Gieq�(�xfZ�8��ˠE��w?�a��0�������/�������C������xV���X���R)oeH�D���>�7�D�ĿI �f�������B�P�_��kte����
(��M ˰���#<ѵO���Ȉ)
~ix��7�]�]��a=�p��������ֶ8�wx��r���QGy���/S��	eh���TR�_���,��@��@�u��31a��~Y}���'p�w�^�����`C3ޕ�~gL�swt�%5�H3gۦ"��2����܎G��.�|��?�.��`�/�A,I[�z�4��eʯ1�+�s����8WY�Ɵ���IE������	�i��+�R��p�6y���N�Ǌ97�Šo9����!<I4bsrA��+h]k:
��5K��J�L�S����:�y|�PF���O?�mɓ�X����_�'���yY�/�mG*� ���$�d�T�p��d4��?(�%�nx,��)�+)� �o�G��d�F�E����;��[�*#���s�L�~.�%���lu}eBr3�>�t�n�h�z�pt��Ȧb�vK8N�`�2<��F��3���eƺK�d�te����6?�س����{�G�7��e i��x�r��椄��Q��$(��P�}>IS���%�'����� 	A��Ί'R�q��3G�`϶5N�bHT"�	��PWJ��A�/�RM��G����EN������
ZX�X�^�i�_ڒ��`�s�\U� ��Dg����B���3�&��&�0�+c�v��\BQ�v�`|���Y3�_�4�ܴ:�s��]��/��iǀ���|^瀚���)p3�!����_�T����_��_2Pל��z�+��?A�_�����s���1j@��?~�e}!j�B�GG��$��?Ww�O���i����E:������6}�:�ԔRO�޺����ڰY$Q�8W͘)���J;s��٢��SCr��z�h*G��@��������V����{q�j�.,��ڤ��࠺G*�j���[�>��ͭ,�V��&#��C����)�;Cھ�OteJ[���D�C�#�#I�LD~����������w���Sh���ƛ���d]kh��
�׈���F�֫�5:?���&�4���&�E�ѕ���W�]1g�hҢ���}�-�(3�#�kلL��`H�U�ss$��yh6�j��[J�~ֵ	9V�[���f�O�'�O��K���eX��Z.��ҒJn�_ɤ��aF�8C��M��@��4� �n���7��}]�]����$4S;h����Eú��]�5��_JF+�90��r�:r�͚:���s�Ṕ�T���
�l�j��}v2�ݻK����\3 9"4�u�ɝ�\:E~s$Ƨ�}P�>��K]�������2�,�+̻�a�S�ow�rG$O[^q��_0�t�|��k��ނ���'1w�'�row��H:�f{M�U:W�ƅ�"'w�;H�֜���7vp�mR�S%bg�y���J�;�rJ�y�'��6&�]�:�{�ѧi��{D��azU�Z �yb�ۃ�:����'C�[�8~ћv�Unx�Nϣ۠c��_w��s�=/��r
7���gs.����PMfQ��#��)�FP�)�;
�(D��4�HE�A:""-(ꠔP(]�H'�z �$�������]�w_����Y�q��s�>���v���\lUu��n����p�e��^�i�kWJn�b��4-��/z:����{�y���hK���q&�j��|�{G����e@5���mR���ni�q"n?~pb+��cV
4��� ���58�w�����Tg�ON�-@nn�Ȕpt�hB2�>Ι��^�m�c:���f��n�x kr��6��M��{��n.���]��	�^��;����w4������(����?�D��O�?�D��O����Q,w�}��t��������G*�a�j��8��ess3������.S>�.�6��E �M5;ח�fw��<G}����
,�KD�r�䕏(V�M]wi:��Qz˽�w�ƈ[��N�}�<��HS��ȃ$�Ra����
@:e�I.����x���pj��E.����͔p�4(ES,w�5>5S���_��Q��թ.��:�q�d����*�]�O��_���(��.��k��B=�!���|U��5B(��t�X���n9,�U�P�0��f�O���Fn��g�WW%����{��}n����W¹��~��O�
K�����=>����V^<�${�n�۷o��~5�T�P��RI-��um���dP��k��9c�4qM�;y��^H�/^��@��gyp��2��Í�Ύ��ן����.���<��}a��dT�_�)/]�F�r��)D��oom�ඬBH��<QUES ��HҾ���k �=��q����;Z��j�[m�;F�����	e�=��%-�g��V@yG��*�_�П"���'��FH	���\�t�α�[�Ł�2���<K���w���~���'kO�	��Úl�p������Y{T��2tJ���H������\$!g�7v���1�����#�#45��^��@�!�j�5ߏ�Z��A��0z�֤�hȔ`��LW����`���!Ͽ�0O��No0�65���]L��X�ʽ�&?���ի��mi�j�,� ޣ���D�%ni�H�!��r�cD�`4)A�љ�<��n�����3�a7l��(pUY��u�8��"qi9��bBi;m���IF֖�J�?�)�:�G�G�r ��sjϏ.�˯΅���\��2A�i� �咱��&�=����DG���1��_�V�yɸh�;�<D�x��y����It�����0�#��xM,_D�*t)�f�K7op}�%�q���a����m:6|
��1
����
�?z��Z���!G��l�y��,��b+><q���@\}D /}��~4���1:\ӟ�}��h��?rZ)��u��4g�����u)Z_M�zN��; �E~>-qͪ0�>u^X�M�M���Z�l�%&�ż^[��lME�Ѫ��PNvRMJ#�F*[ :#'Kp�?��yq���l��g���$4�1�fu̪��*������N����T�ՠ�'�k���u2�د����[#����jl6��p��+���u�ܕ�A��Q��oȺ���E��L�����?o��JQ�BQ�ZG�
�[�UK�]S��#2���H�����x<�.�8�5d]��{���
�zN
�覻o�����\*0pjE�}�@v��}c R?W��w-�p��v��8pbǥ�};�����������_��y�����/�<k��!��`-���Y�l��dԗT�������{�\�דN׾���6Ɂ����YJ�vk?>HG��sg �0yQn��k�4F$�5Į�b�Gx��U u$H�>�]�k��`�<�c�b/o�D]�^�����7f���������1?(|�:�N2����1��wא��{'جn4��>R�:��#�<f���L*|ϒ5�x@V��Q�k/%4�
�
�uF���'�$��n��A缢zE$T���������f�\C|���P�Θ��#��RY��819���I�<���o��C�XǼAZh��+���Lq��M#,�X�8N� �4p&N}}������-�m��c��+X{A�������>�=�F-����kLh3��X!�����m{�p�{jf���c�����y�BE�f�#E\L�L����+K-Ǝ,< {n�0�Cz;��\y�L����M��2�����:����Ck��}N����������TmJ��h����u�W6���߻܈���1��E{qa��X�z�*35�	 � ��C���}��E�jʜ7�z�LhC"���kGN?�x�&'��+�C��ܷq�/`���
�������y�J�W�@��EB�_�#�&S�����?����
�1F����ӉK����"�&8�S�[uB�b
�T�2C]+�I��ty����,��@�x,@̺��7.5v�/��>* �/%.�>�V�^w�J�#�x)�����S%[|�/��;�o~� ?.�,��&>|�l3��t���Y��������w*�=E���� #��sI�ƽ��FD)9�k�B:���IS�ݻB�]C�W6��;�_����x��r��y+�I�0���ɩ���o���|Ȑ�F�]��
գp,��Yn�u2r�ע�à����K����z��R�,�tEҾ)����{��؍���6�X� �G�G1um%$L��I�j����e�0�X[Kv~�>��w:p�z���ar���p=�L2:��ݶ�풏X�d�q���]�#*\.�#�ݪ�+_+�2�30�r�j�������<G.�~���
oBյ�]+Ei�׶2:�z�!y�P�����k��]���t�A�TI�����\)o�{@\�F~����2��_�k�^%��(v�_�n|�-O���H�Mhs�z��Iv��}q�k ���mÞ�	�]���@�؛����,�w�Q�qKaa��X*�R��<:�J�S�`�W�iK���B	�C9�,��������D��'� h�o�TI!/X���M���5z�ڷ�/�Y�qĕ��\�C^�����������ג��$S�ʹ3ل#V��r�O�ؖ�p�w�f�t��}W��S�\�+�7\�N5���f�]�p�"[T�D��ۏ�_��uvv�f������_�.���{�a���W����>�5�"�KZ~���J��\S����^�zspГtGW�� 7;�#xq��7XM� �i��D�F��u+�{��|����[����{��Pp��J�����Z�?��=���4)���a�hz��GD	?ݺP��	-�VO/d*wM@M����
<fBU����eW�IYɺC�1u��S��������5���H�X2y�5V�@޾�+�. l�5�aeƄ[n5aM4�Ɠo���S�q����|�ˉ
�(Ș�����K�Ԉ��� ���/�	�v�+bkF�Q��#?*�Ԟ��vШ�~��|�����xA��R�~�T�^/oQ�0e�����Ƹ��������\�91��A�No��?�bR?]Į��)&&�%���e�U��ѽ��3�2���$�}1�DQ���[��6Å3!	9�o�6�?x�T��G��e`�Y�-+,999_�\G�͕"��.���܁\ȷ�X���\���Jy������Gp��L_;��y88�䎳 n�����*K[��+/S�_���3n�)�K��H�[���?r���u�#���<V�k��s���2�(����B�Vl4U��dqa�3�
f��ʄ�X�$;�',�����yxr�RdY�54�D�>����ׄ����O4ϑ�m�G��"��ɗ���P��}C�Q��sؔ¹
l����A��'ob�pw�>A�q�7��{�8
�hi���8A���=�d���~���$�Y6̄Y���e�^0g��}�-�˸R�ޑ��m	���8g�4�ח�ó�h�3������>7��>�o�9CS��5T�j繐G�B��\�3ԝ�����`�}M�e#�.�vK���*�]�������u8>F������e]ԿC��u�O�L4�.��H�*�nޠE{�F�uӏ�E2W�
/�+X�	R]��K�)�B���W����u�?����7�ӝqoI<��v{�e+�'�x�VU��{�h����=��:�eQWV��R�bg��vѾ�Uh'�n-\�Q�/m�
���&]f*P����8.(�����d��:3��	!��â�;����7X��>r�~Tu�=gb�Z-�>_�["H�n/�a���K�{<`��,:o�;��ci�V`�,�h*�i�XU�g���^�T�bsr(V�D�����U�_p���K��ÂABe����f�:���q�?�V@��RQ�L`na�ix@�Z��ܞ�����g���.Kp����Eb����]+kd�vz�����,�>�;�I����p,��Ç���]k%��$Q}}}���:�5��9�E�������r���Q�t-{䉵d��x0���>x�<K��3v�����0��m�� �����y��䃔��&뢗�'�����i~F9!�UH	4�Cu�1�� g�濖�L��؁��Xy�r�\a�V�Llnn���t��S�N�-l���'hӷ
�� �;���/����!����_�	N
F�zf�����dt�cFA5���^�UfA�Zu�9)i�lA�d���WTo�	z$ ��F��P���n��|�����B`�N����G�Xg�dLyy"�>�wB��߇��\PX�)z���2kH�E��Ӧ�;��#�:���t}�6����5��Kd�����}��X�L`��.��~��P��&=NPY�N�n�,��/�|���S/��g�/ʮ�vyX���]{b�滆��3T�d=<�$�Xr?��CF����gryX�ԙ��i�����*��0��e��\;"�ps;j�jr}Hr��%�6����x�P@����i��=�]��pK[��[J2�R> 0�7�BKl�/��/
�K_��	��t��C�LNNc�c���q��=Q�󆼞��^0��Oy��Vg������ e�^,N�����d����.+j/h�Nq�6�U�&���Z�fbr���`�>�&��lsFe9�X����[����5)����Q#�|h̢+� z=i���3.Z�<11QǔȨ?�4�� me�p�IS��
S���Y ��".`��ԙ��\��ҏv��_l\\���n<;P�Ԕ-�Mt٠S��(�������շ���`N͆�_������q#F%4?�:UFU������rz�]���~��\�[M�n�g���>`�S[[[��;�����Ph�67w��7�39�-���
���CX�3��yh�R��j��H�tvvf�'��X4�<`Jj����H�?�+F����^;pr�����e�I�+<]+ �	�zzzZh�t�B]���@�%SiQY`ٲN�\��R&'ݔ?h����:]�V� mu٢�f�&sh)�fK{�=<��P��-ҐM���N�@�~s�5����qxju�K��h��lv�2L�Y�ͨC���{�3��
9��S ��(�7���_�+oI%�b**-�X��(ⶵ٩I�#\e��d��u�(]PQQ���KNO�+@00�Ծd��|�UN��DGGG��V��.�����)���n�,Z��e�nL|�tG�e��fuH�����8���>`)\�کEq�F�E?�����Ō��f��i��"_���(5��׆<M�u��b�B3���<�C�j}�x���އM,��:r/YF�\"��"E���=�v����|b����R�=�W�ta�޶�璋7z[��~�y�Zٛ=H�^�C�o��)��s���=3]���_w$�;o2p�8������wށ8����GyR;@���v�ꏷ�99�������/�Uȳ��>������y222+3]=��'`���*�����CCC��&�}��:wy�?���9���������_h��K��P6��&ݴ��ٓ��̃��%c{�K"4�Z���4�~	B&���1rUN�h�td�#�GPs�MH�3�%�Lm�jӛcb ��q�t�����c��;��]�WٵJDPWV�+��.J=Ӆ?Z��N�3; �#��!��1N��iN+�TZ@����B�vu�-7������k����p�?�꯯�N��y���V���o�w����bS:7��Im�����M��D�����a�����_OA?*�<;��>�f�_��'?I�x;9�Ư��S�c�Ϝ�{7E����W\��h�	xv��ġ]��rq)Ĥ�9��t�`3G"E��$�����S�!�>�D	�%�B��|]sՇ�<����K���"���k���p1���� ��vK.v~�D���G�OS�ͪ��瑧��9�iԖ�Vw�,,縕Y���r������!o<_	õ<����+��������n�D��7�_#���NC��V��i��|�n�m��˜�6q�&����P���Ē�.�B9�����΋@7�!T}��ƊCW��Z8�۰�&F��b���\���e/�;���0a�6&$�"]\\ ��(,\H�K2Щ=K4��w%����&�%ʆ�25I.�;��U���#=�VB��°�F�^�ТT�"$�z:�5�:$N�8۝�a.��i�n�C�u��!��5���bJdVݥU%R[���s-���}��\6�	��!�����՟�yR��?_5��r'�"W����=�:İ��򻰨�/[��g��ot3�55R|!����4%u����r�����`sV�>�p'�Oۀ��M�ŵ�!"�8w\1`�<�*������g��W#�^(�k*T������}q�%��w*����*ɸ�[�Vi"J����ݔ�aQ��0Y���ɧ�a�E]��Ο���	I7�:�����ܣ�G�(�[_6Z����X�{j��y˗�g�Z�U��cw�:�1�%VI�G4:�p�
�vy���ĕ
+;��0i�_��Z����6�M�ǒ�
/�<��@;�DݶBM�U_ Z��՚Ҳ]�>�2�amu=!;��1�g����/5'�ͅ��"=�s�k���v*���G�c����9�<��?��O��s�d���m-���}zG�e��02R�R��}�*��_��5q4y5aC���G4��R����e���W̌����������#oF0����~��Y��@�~�P�vrPk�V�q����|
ћCB�~Jh��GO�r��-u�PIԅ��K����ِv�Z<�ʚZ��M��8E��v'^�48�@���JXc�	�<2"d+�c�����ҹ�4�$�{W��z���>}hY��R%��5��~�q�h�Q���k.�y5
��wv�W�g����ɗ�%+]"X����.��MW���R��3vp��t��ދ���T1x5Z�h�n]u>D4�צJ�ۇΎ+*T��\9���}���i����|�|����(^���s#Z�5�]�vэ���ĵT�Q��]���-�JL�/u|q��dKn�bΌ=Ito�j�S/k���E�^Ws�:�)������UEBN<��R��z}�å)�҅��i�7�U��o�opq�q��e��=9�NC���mP��o�󸈫0#׮È�O� �y��+�ֱ�/SF9���c}!ޯMרH�`�բ
9g���(�Ό������K�M�|q��w� Vr��$����8i��ܝ�;��W��!���@#~^���
ǖ_2Y�C�7H��d���uk�B��X��,ת��{�l�K�W)k�mPͧl%��bdi����ң�LPDs/GӪ�t�m���m����XH�v]�&����wS��?7, �=�Y�пw�/��W'°K�J>V��>t���O�	Q	��+��oP��l�Ǘʩ.�f^�(_ݒ��͂۴���9�}	��{�*��1ۧ$�g"���XW����Cj���9*T1a�T�]sv(	g��R�¼h��-\�yA~</GfKO\N�y��O�0����%�cɆ0�A���Z�����G|��4 �Q�W���q�������=y��e�zf�I�\L^jG��\B�Y( /�{�J�w,���	o�'���t��g��j�M��MT���m'g*Qs�6>��"�ǈ�xo��:����sTH�W�l$�{P9w�[�U�Mc6�of�Q�𴮾�Qu������_0c��+�/V�����[�9���l��G��5z*nI4ή���l�<?3��5'��:�n���&�B*��e)�	}�#���Zm��WI^i�a��-�+�o��U.仰�u~�;?ZC���Ĥ��l�
�D��#L`{�s�7Ҫ�b�}(�4^k �l�'[�l��\h��$-Qo2��T6��oe�����+����z�������@X��-�8�]�i�\z��`x�3^#�]Oh�u��Ls�r��X����V�#�w���׈�\]e�H8��QMu�c55dlQ�㫧��)�V�p��2k���X_���xZ�o#n�M�Br%�$�ƭj�V�/���r���N��&�^���mw��*/����M�x�c�cx���������7ڙ���.9������a�k�H�å9/�#p�7&ν�c������h�	o��PO��S!�҇Mn1�B�8W�RH���K>�_�Q�=�׍��Z;#���g%�G��l^)V,����-��yiɳ`N���Bn!G}���15/qCy=&���4�����dM������	�{R�f��Mѫ|���u�t �`���OA�9�wh�P��8.�g��{��h͗���Xʩ~(9��*�u`I�r	YTekd�qA�4Ds����ͬ���	�=�nհ���� 7�{���BU��B�����w|�gA�:��D�l#��t��CIw��ê#����β��Ȋ�e��RM���v�q�gc��c4�3s��^��b���h��n\X�@�5&��F�/�5�����S���ޭ��f������=xr��[���w�i�8��61�����!��6�%'_�kظ9	kT���;���plX8F?Y���9��Ԫ���P���)1{��� ^�YSs�B���2>Y�󎭭�y)-P瑘�m�vcU�c��G�x�����<�q���޺T�5I���Q1N������;����k"q�.#�zzzK"���YQtC7�4ٜsaxm�X��Ƌ�J*��|0Io�F+WԻ���z4_b\�����FH��f��������@1��:��j$Y�.��+�!+���c��ѹ7A��!5,AK_]�\�_1�0!�Zc�q
1X[�#�&�sL�^`Z���)kw�E�W&ʀ�WY��h����,����%����j$�ZV��x�$Er1����.���[#ۄ|�(��p�Y%a��Z��DZ�g,`�q�ڧ��.���^t#�m��'\�4�<�e�
4�<ahZr�
ȝzz�]9�)S,c�(F������H�<�-9hX�aA��#��lT���oe:Z ���9)o��f
X��լ��W9y�^=w!����%�O��G-��8L�����ۡ���-�p_�3HC�� �)5v���9�CV�+ҽ[�������2�S�u�QUz=�x^R�Sc�O�	C��u��~@$�ߕ9���<�?�R�1�	4�d����8x>�Cn�xn��l�xt�7�X�#ӷ���Q�Iŷ�ͨ~mw�ʍ;��ӡe� ����_�8C,���$�4(�V'2�8�hiZ�ϔ��� ����]�Xl���[4j�>��]�hğ�,'Ʒ���3E�+X��ي��uu��k%���T�;*�%��#T6A��NC�߰��kZX��\j���NL0��`r���Ṃ��'�@�d�����\�Z��r�v��%o��s6�g=���K�$,�ñ oБ��cG���[�l�<�#x�y\�(��[��j�YR�b������m�@B֭釋0�z�e�j����ܱ������)�f���c-�<l,Fs$b��7����69)�	�ל�3�7�1�T`��]�.{_h>yQG�2���Y��y��.��쒳��#�|/K�]�cā<����y��
y�~�4i(�@bg7�rYG��N�r�զ�e�<��E^�䜈J�=6��E�o&b���C�[_���l�a+��?+��d���v)�r��k� a9=�Q�
t$"��	y���5�g'�ȘU�ѵ���0.����f�eǎ����o'?C1�.j�o�
T�4켒e�� \����3ɍ��4ߚۯ0�����=�Z~�ϣ�J�0���A�E��Z,�F[�P�AU�؁��*;�P[�Tp�����٭C���)��������Kx�\�ĭ��܋\L��9��ҷ��{�Q\�ّ8��;�Y��<��T+�a�ǛҷP����I5`��������A���v��کk/��o_��Ӹ݃�|T�(ˋ�.�'���ߏO�\#�����{���/!�`��{�a=I���KA��r5]"��.�FJƥ����B~���U��Zv�Z»�\�8w ���U���9<h���c��ނ�ԓlmF����	Une�������W�@!�kڂ_h ي�ra���03/��w�����{��U� D��rg9�D�~2x%��������@<��T.�g�%�/L����4�`��S_-��^.T���ު �9b�8��� �����tՙ�z|�A��*r�4u�7g�Z�36�7Ns�]f/KK�X����2i�o �xy�d��0[���Q�����L$Y�JG+i��EP��9t=���r�k,޻�2'�9݋9�W]ϧ�`��F�e�/�:a��z�a��Y��w��5#��6���O��X|6��=���θ
�@��Rt�W6р ��Pէ���٘-f�����bV��Ǐ��ܤ��
�ζȖh��I%��#����*�PY��6����X$%�{��,����R��C��`zV�G�b�:�1X}۞�~5�4)XSs�]~� �|��k6D��,��R�Hҡ΄Zua�@�D��amHUE�9��?��A:�*�hQF����^�a�����@X��_f�z7a�k����ـ����d��D �#�h+��0;+y�tLP��֜��������0���.�w����m�m��}@�>���ʒ�wu�Z1����.�[�W(�l<���?39��R�j�{���Jl�����m��׉�%BCbZ�AM����D��bS�*�u�z�V�q�5MBoRԕ�,{i}ix���İ���~��'┋Ͼ��<���k }�j�Y��WGA7�݋mN��?�M�B���[Z5!�4��^���9���`ԣt3������0�z���a@��P\��bsG�����ʂ�k��H��<٢����`xu���|�Q�R�՞Ae<=3R�&�l�G���}Z�j�M	��d�@�"��Ճ�CE��#��4ݮYH�K�T��zh�[�J����(�p���7R����*��m� ��17M�Z�H�2am�O�����1bq�$mc:G�Ve�sd��."L�G$UWc�5��4��!lY�Ӆx|)� )-�<|��ǝ3"Q���C��[��Lu�B7�6��a5��Nꌊ��J���a�4�3�uQ��bQ�yM�e�����f�95u+�x�����h[Ȝ��㒪��5ԵӶ[�Z'������L� 4)j�w��T�J`������1�2£��uO��Uq�-T���Пcgq�;LR^FA]P�ܝ�Ea���[7��_L̟\hԲ?_m��c��EGPO��)�h/�*?�GF=��6 �ҡ��ߪg�y''?��]6��ز��73���*"�����1+_O�(���^�i逭���/�h-)7�(+�����+;PR�.���Ц�����7m�^~���q�7y�j��X��G��!����?��M��vJ�4���wu4��C�j��2� ��>t��7Q^@Yʻ�ӡi|��v;��>J��u�OQ3��5sV�Z [��j���P(����
br��ۮ_`��vKX�C.�Dc�gC@r$�IK���܊��D i�ޏl��>�@u��"i�/`�k�qg�d2��n�G�j�5�(vv����C,P����Q�@�5��	F�7�k��Ҩ�v�A�?X�vg���/�U� -_Mwܑ�7��op�����@��u��	M�.���<�ܫ���5�)���F�NL	 	�(�F˂�2�q�G�W�4����0F'48���H�`5��V��YTl��[���Tax!Ǥ�)�����R��(���?RQ`�>�q�`�a纼��]��.�՚�p

��J����l�����+��/\�Ҿ����L��Wy��H��Z�R�������J��ƨ������v�+�[8U�V�Q��)/!=�5ש��N��;ŧ���zm.�L�oB�Ӊ+�f�����A�l�,��3�i��ã#��WR�>I�3 ���9�$�h͈��O��j��VZhC����^~U���U����ZH�R�3曄'V:�iW��}&�Y��Y�^,�,��ʓw��
l�L����G,�l�	�1bN��&X���kX.�?$x�@b�%P%]�TO1�����P�ˢM�k!���[�^|�;<�I�h�>p��͛�;�U�RKv6�ޗMO��yj���%�K�.cP��k���
���X��]u@P%���c��`�P�%^ JH_�N/�f%�i�q��Q��,O�q������+Xь7�/}��3A���iɕGF�}F����S��u��rer�$y05E���kt�'MF0���l�F�N�v�p5�l���.0��:֬�S�霐�ˍbz[��bH�E|�^	�c]�,P�3����6:��R�ԟ&=��ZF�5UC<�֯_��6�Ar>}u�-��1Jڇ|�㿖�k�Ԣ��ÏT[}��&����4�&��yR�;}ݨ��*�Z[�e�!<i�+P�P��^*Zhw�.����[�f�M�識�1A��r���O���T�r8Y}�ՏP
k`�@.��q��z�U��(f�'�/y��<�_���N E @i����J�אռ����K��H0�m��x�����5#t6�L�
V�淐����8Uc
�8/�	X�.1��h�%4�Eh���v=����g��2�6�Թ�q��=L��j�FOC��4��N�Gծ@I@�@`@]ZI�@g�ݾ�.�R�F!շ��V�=!�#@�^tC�����ٍM:����By��$�O��(4h�n�"F�M��N�M���lm�[E��z�:��%��}Y/��ش���9���R�H���gh�!�t�w��8�D�fc�w�q�hrv}���8�Tt�q��>��V�S�>S+�k�	�Mvx�7֥`�Ɉቘ������Q��U(�!�I6[��]��c5��_�ʷj��j��+-�ǫ��9�.>�幒��s�0�YB�JU/�K<�ڄ^{{����(���Z���4����P�M��\�`6�OU�R#�.�+����©�c�%WS����,K	�m�C���L��U+*	4�O�Z?�|�8��_w�
��+��\aD�I	A��������ܒ��|u�E~?-�Z�Bu�6�A\������H �/#s �W�ďjjO�x�vO��k��7���4�	���C��ayD�6���Y�d�����'Y9���q'p��z��B�i~���S�g�33�x�T��%���{'�!j� �O
��9�4�l�B���Q��V�w0�`���Y��eM��٨g����Қ�Q��'������^g����Åѣj��K�=��j�#HS�����"�!�+�;�N�`W�U���Ĉ��D'���-�r	@�ԓD��gG�B�\yWԳ�t\����s��~cE���'*3!ސ��4�pѤG1�8u�^���P���!��e�e�k�a�9���þ��l�~.Б��zFZ��T]i��+��τ�|�
�R�I2alY�_�'��?$1 dI�92n|VVǨ��-W�L�p�TT�)<��xT���]�bƆ.�B�JHN)We���{�%򬩥�i>^П�E�a_�Ɖ,�Bi`%��ƨ��U^}S���oT_�{��7�J���-Z3��{}�CYAt~!|��Ja��`y�`�R`�S��]3s�$�(��֯_>�6
!Tױ5aa��1�4ػ'g� �t�_̛�=�����v�u����v����gl@����1��*����ꗆ�M��0�[-�lxA;\���`ݼ����1�|p:H�]5��y���yŚ`��GkLô�a���O��m�k����13JқC�Z0G��RG��e��������D%Y� �77���gxAmWk�!���/����g�s�b��8W�|FY��7�%b���
����X%u��>,�֍�_&:�7R$��zt񵒊
g|�u�=䒾/=G���������Wm	��=�ԾR���RB/%;�d$�r��s��JO,���澄��ڥ������;F�`v�������/t�j��+�a����{���_\������_�����g������V�Ż�7PK   6f�X�;�К> � /   images/277be1dd-7489-4b2a-8eff-ec6391927629.png�{�;���w�t�QI��PI�T��pʾ�{ن�M��T�,!{ɾ�ef����1�a�ӌ���ܣ���{���\�_�뺺�ܟ{y�������D�s�=v��!M�C��Q���{����q��o�4M���G��ߏzkX�:������VWc�x�O������n��t��t���:�{;���qɤ)�:t鐦�}�'o����&�;צ�p熏F��_�6rgLT��I�.<����6���L$�<ʋ8�j�1^���ߗ�
��{����ޔG�'DD��fN�Hn`�3ȶ\g���Y��W�SO������/��X����������l�[�$��6>|����}9�������7���~����?"����#������2y�g�L)j��b)���_��8�n������]n����H-�opm�Z�`����}Qq��S����'{�2
�X�|��Q���wx�yx����̿k��ט�Иy%�*u:���QRR�g���A+pƛ��L��A�ĆqUk0��V�c����c@�9��i-b�xo�Q���Xj�RNB[?��ayyG-(H��G���{(��HE�A��iDU̐�~�CUT)�\D�ōJ�L����ߢ�c���?$q\lXZ��a̙-Mv�D���==y�����Î�J���(�[��73���Q�gS��q8�F�n�HxN�"sRT^^��U�LLɻu���z�>�M��)z\lf�R?�yY�%�>�z�:�}y�m����I^�������j��beu�V���{!nY�k�PI�����id��q�9!������ؕ�Fۭ[����[*y���w��z��v[����J.�sF�붞�Q�����Bjh���ۙ�z��e���
4k���u0[���	uXJ�a�C��cN���AOPvXRhw˫ciSSͺayY����ؖ�˹�i�V~���T����no�|������9�{y73�ԩ,B��F����vB�0��!^���;/��G����{�t���q�Nk��rr\���v�)��<��p�oUCl�`c�!��;�e�] m����eC�
@/%r��볉V��}��>E	*I~�j����g7_���F�g�%�=���{�C\Rλ|��}w�'�"
rN�v���E�)� a�:�c+�����9�R���F
���6������+�c�����i�};̿���Fh�.*���L��ѧ�����wj��dk}i��A�9�~�~}y�=\B_�]!�⌟揖ɺ������eeGq�7�W���v�RU�ii�jQh��q���U�
��`�ID� �˳/s~��V�~e��`K?�@��J̮&vw}QO�gU�O!�k�'�&�ؕ�����{Y�D7%���1�0��� �͘8��/�m��4��#,�<�p�Zh���m����(S>]j��ߗ{�ӵ���YH��?���FB��B�?�UT4�n��+�v�idd�������>K9G����M[�����y���������o�֥�F�U����n&��au�g]���~��� �m�cnB�`G��y&i�E*2���V�j��mHL[���ꮩ49B4��"a[��G��)U�X��v�<�i��<��f��3�A�Y{��q�Yv}bt�c��Z��}l�O�[���[7|��9���hJ>��D�"���>J������@�/��].y$@�4l�%Ի�M`�|�1�R�i���R�?�A\�V��ӕ^��~��7�w��]L��p0NJPg�y�X�LJf���&�e$ܑ�'�7�/��)��m��S��GŞQ���-8�]�O�h�ߚ����8X�e�jK#�^Qь������Y����5LK��x��ڹm���$�ቷږ])��7�s^M�R�ep���a�0<�퐷KoT�W�u����
pl��`!�g�@}&�S��C��Q���1�')A��=Ć��[VvD���s�M���얩%.v��ŭ���иcc��m�ـ��w��B����dG,���6�[�a/(R�
�HIj}G�[�?Ѹ�T;�`��`�r�rq������B�)l����*�����)���q
/Q"�>ջWQ���Cwe%Ey
�1�I�؜��0�b@^��|�$���>� ��a���7�>�-m��_bF�<��������g���X�R����*��C�h�S�oiSJA)�O5�$��q_ٺ�b4�h x�ʎ�r���A_��«�hV����w<�8R���@ܼ�_�Im�����hKk��ߠ,��d�>k��?��S
�S�,��ᒾ��y]�`&��@�t�K�@N��KL����䞄w�z���cbc��n ��S��?�ׁl.��z[�={������A����<�;�+ai�6%;t�j��N�����?x@����sG0hw��$�&f�<bbc���+:,��!�j�ǌ�����[R~*5�a5���WӅ�C`�FV::�N�6���d���船�Ɓ��\tNur������]|�2ڍ,Q��c��D,H.����W����N+O[>u9yez��������^��M?�\��1^�W�c�x�2n}�[�^m��)��}�-_	��M��+�x�7�*A3zz�X��S|�5~� ��ʿ�E�@q���;�����Ǎ�I��sr >؆�����VI�d�z����ܯK!�lV���5F׮���//?y`��Ɣqrq���\P)�ٟ��54B��_�Qkc3�{��z��_$d�}�W�S=".�1N�𙖝Q�A���P�� �����7�4�xaX��'������>9�Q?l<hW��'��|���g�f����^$$p��#�w7�)@�g��#2���H`ؿ	�#m|n�ꞿ�;�jF ����H�q�@]_��<1nC��SOb���P�
�J�� mV�xꊫ�v�ʃ�j�X]ի�~JL���$�HTdI������y�r��d$�3��b����/_��<�\�3�+f���-HW����Vh�7��
ţ4m��������V�#x����E�߸^�K,���1`Ja^�a�j��V�ab%��n��۹oѭ���7{1� ޻/��������5�xt=ca����,OX1 T/���+<����F�OLI)���'x�ʿɎ�Лۈ��I�tP�ٱ\�2��׊D�A� m��������E~#�k�zw�tV`2���Xejv�h-�k���\�a�QL��O���sFv�j��O�����5�֖����Ic�Y�f�yJ��f�h�n���+ڍ��B�хFl���m������fڛ���f$�{�p��� �C�C.����mЖ���	��_�l-�j�9�>dPDJ���Pϒ���nVf(�"N��A���;Q����W]�Wø�]����!ƅ,�o����.��.O9��i�d;L�,���)]�Q#�y��]��K �*uR$z�AAʈ�q��c#s x�qAA.'�G���-�,�o�����������<�B���ߕǶ��|��ez�P�V6���Y��Kn�
�t�s�uF}K����I�1"!��㌠X���ܠ1��W���н_s�����+e�ew�C���]Y�d����(��Y��O�io��Hp�*��������R�����A)(R�$��844��{C�������S�Py�5Zj��ޤy��H���yD�Wdg-H�2�]�y���j���>��0���*�W�A"�'0>��jϡ��r1����A+�#Ϻ�ǔ_����ָ��'t����I�
	k�N��C��md-ZP��8�Þ���K�C�MWة���v�6gQ�# ����`�� �C}^.���S�.��3�k	F��Q2x��E���K`Ѕ�g��XQ�m��e����㯵`_N��d=r��,9 8����gմl"�^���ߟ\̔qB���� J�UH�
�c醽��:��֧؟B�p!v@+~��I����'��7�P$Jb��(���>TJ�;1� >H��c��:����TB�V���͛���(�
�ߠB����a����(#�~����Eg�H��D� ��'� f���]���Y1��x�k�$ r$p0+�#�/B��r�T'��B���,XvJ�+H�f���U��E�W��
�&c�f��� ��v�z�D�aP�\�\���Io���M�^��F>2gg��F��A��S0�PP���Ǘ���򙦬P������")�]�ƇՍ���g�2`���	�A�-�XR䅊Ա����4%��{�K_9��Q��65�s>��S�+ː�X�dUhQ(f;|�c���[�{W�#uڿ�h-�:��,����80D忧�I�"0�a��I��&`ď�[+�/��@��������f����F�ݏ#26��X� ��N-�����O	}���1���%u�I��|�3�t���#�"��ĸ�-�=ok����~�
�X�3^47�a�J�*r�0��c�uKZ�Y��+�a�X�T�]\�5�� }F:���D;X@��+d��^%�)*2� v-3ϑ� ���HA��lBH�����>�@��u4������{\hʠ�Q5�4a�_��?��al���ķۨXk@��5���>�!J4��\
�icipҿ�l�i��`.��?DY�my�JX)W]|���Fc����"U�r�%�ս�r��A�֪���n/�wF����A�6�^* ��?�\����C&h�A9���0o*����p��<K��� �>7\$���(���zy6�����E+���.�;� I2�!�²�j��`?�V�,�5��5��TO_���$n3ǥ�l���������%A:�M���iD�@Ѓ �-��{���;tO�������Q�H��>�*�����HKI��#\z�x|�7�����{��w��CVK
f����h�i��ݏ&"��aJ�/̾��?��D�<�c�p�6�.ض�>'����*�	`��e�|�8?�G|qBb��}�H���eL���(Y�m6�FB��3�V ̽��z�y�c#��$6�pF;��"�g�]�ܱʉ��~F���%�������-,��*R�S
9�2W��|��o�Wxlx
�S9�۩���
Yw�L�Ĕiщ�#��pϹ
��ŸF;�����<0`��e�b�|Kn�.Ku8�x���}��֗n�A]P<�}�&d:b	Ҡ���UT{���L��X!==O�Ck��HE��̝�^@2�m��gan���$&�����6�����l��48���՛+��$ �O�I/	 ��	���<G�V��Y���z�I��細������&VVP�k���v�%}���5���,��C��L�?c�t�(Փ!?Y_���Z2��TI�֤�ʾP������gU��Yw�k���Yh[������F�S���N�kM�Zn����k6^��r�r���a�����{�B�ю����ej�,@ҳ�S �&�u�_�p��Y(<����?��;~qO��3aH�<��2�2����6�s�-É�唉�G�\u�`�+��9	F��e�/e@j�'i� ��b�����{_����8re���O%�&���Tk3��c�څ3f���_O��������\�dK/����;��q�"��8���D8�Q�	Y��u}�%�x����
/����̥�-��}9�������!q�s�)�B0:O<>)�����5��"�7^�5�u�Y�#�:)�.�T�!S/�Q�B;X g���m�lG���b���M�#2��Yo�дW,7���Q��!�
��*h�����E�V[I���^�!s�y]"�>�����T]k�턻���o�C��{:�J� �7xc�w�rFz%B�z���`N�A �OBc��\����[b��3�엤oW�'2��_�w1������n�V���jt*�yn�s�'�Ge����L��j�ϳ?m7=����s��e�Yav�Z�?5ۋ�<��̫&�V�nj���o��E#=F$�|�*`,<�ʩ��S�
@�C� %�:�b�;�  L�6R)M���Ky�qEN6T6-'tl�����!J�<��i��[_�e�ͨ:�?�������Qi�J��
�g�=�$��~*HJ�X%�&�>��%�k���vQ��o1��K�;�PD�Vx�m���/\<k��n�oZ����s�G_�����/�XU/(���ȟ��y/ɾ�t��q��]~�|�B���,�N�a�נ�f�����q }�e�&s�S�+>*ǘ�B�#��9Gؕv��[w���0���m����:���:�����7�O!���i����K�[5qRR����;Ь3�W:.C���ŀ)W~zw�m���%����Y���Y����ͺ�oP��E:�BL���;�>1�!��9 j#+�ʨ���}�e�u	n��	�9
8Y�4���'V9ì�m�gF�N�1���zK9f�Դ7��=��Z���W{G�@�6��l~�x�
��UzY78.��V�g/g���Wp(��X%��������{M�n��r�1��y��d�n�5�!�z6%��4�LOK���Z�w����S����V��|���94���Ū��'Y}���3+��y�kl�<�]=SQo1 Pf��z�ո�J~����®z0����j�	y-V��H�0`[��<��RS�Ǫg�w�WT��ų�!��mqmw�4��ǉ(p��B��99,�$�ɞ�B	<�fa�w�v'�zI~�~@@�SЍ}���<	�;�6��P�B�З�hM"�A
/͌M`�1��UA�s��?�B����D�VA��$9?	=�C�W[��1x�6�&&�����ܔl\�ל�e�5�f�V�H�:����]XG�P�ǳe�ˋ�kc`<#Y�����$�;��k�u��i�B��!�.�(�Lک�D��k�o�4��� �zʰ'�04l|!0�9�#��#��S��b��f�{�)AJ>��G��6[��a`=emKr���z	�T��@��4�Hb���	��Z��d�j�O���'8ٖ�� ���<�N��+���?�?�i [�X�B��+]��ј�]! _���|�F�N`�� <w.��@m�tG5tRAi�\�I�U%7��S:�8���J�q���.��
�%_�Y���ܴ�(�	������.��.��ҙ��D��ob�Ԋ.�=ٽ3��e Q ��H����'�$(�2���k���B�&dy��Y�x/�:7��/	��#���^z��Ma(���1 �O���B�s^+��!`V�/�kz��l@��)yoJ~��K�-'Y,ch���5q�r��;�V�R(L� ��]���s"�C���GA}_y�� ����-�C���2\ܱ����rk�ǽ�]1	��m�}F.�Q�Q�dJ�����E������&�l;;�Y^,/T�ـœhs�_�D@Qf��g~&��D����/K?�Q��_�9������X[S*�����>���pH�zmT��䝟IPbaL`�����e	�SH��#�B�}9�i�J�"ېyvP�k,11��JJ�Dć�D�9fH�"�&.���k����> )�7fxmH�dV�d�������F�4�����GJ�TJ*��0
��v�>e�B��ɕ��j ��:�q!1�=��봐��@��M��QI�-��*5t���K�߬��״�y`�[6<<�����t$謻���y4�2���7Q��~е�햏�Di��8������	<�-����aLV���݁�Y�����9r���B�#B6g��h����<��	��\�U!������l��Q#0��xw��rx��dk�m��܌,�R	���࢓��5!Hq�Ia0�^i?���"�>;͊��ů�'ݎ��KG߁�ecË��[�l��r2�rNK�W�����l���`��~tĈ>�b'V�ђJ� B����p�{,����Ŝ�K0L�o�AV�;E ��$0�6�G��� Kaw%}߿�[ǋy�$�_�B~\�a2����������7a�[}Y�:��I Ѳ>�mTYr@���R!�߸�:mx.�(�y@@���O���+�ќm�5�r@�����@A�<;u��F�{���$e�B�Hs.�$Z#]ɍ,X<c7��� =��b��E@_� ��.����ėD� ���
��;�IWi1��^P�.�[�.�fBt�m8C����X��y����^�G�6�mtན� }U�;m�}v��u_��u2eW?��6���kk��/�=0w6���<*K�C�w��h|yz��]�-$��=+�7�ɗ䍥��yΒ�E֦^��j�CjK�cN#y
�6�)qƕ�MjfT<�!��޹�2�U%u�6O�tHMt��o�v���tÿ�a��x�!��?���F#��Dݝ��ڿ�v�/�����vX1��Pa_�ʹ��cI2����sP�g:��mI�Kv�6����s\HD��=CZrs�l��=����HE7�w^�>�qFX�NQ�Vb�W����S��N�=�O1��,bX��q�5��,�؏����T����ۤ 4���Z�X��\\8q;s�ۇ,�E#A�F}�k��<�"Q����:�=B��
V�){e�"�;�x��Q�)����y�Q���S!kˠ4}��
 ��VX8����KT����v	 )寄��Ȣ�nN�*�g���'��
Rk����2�*)�N��SK^�cߠ.6G��XO��2O,I���a��3��l�������J$a��J�'�jSݺ�W�iף9٥�^�� ���e��=�s�Ajf�_�Ӂ}�& �~���v6]���d���n�yP��f���6��[��?ޏm��VN���}��Bt�`�P�EFiq��σ���/���h�]�q^Ƕ*ͳ�嗝�?N��n$@����T�$&�1�Z�3e���_���A0�#�x�8�^=�i�)��@<n�(����C���淹���ԕ�� �_Sb��x�� ]��2rZ���϶�	��QEW���Tq������dy� ]/+�9w�6�Ho��lձ�%�9t��6�ݿӀKO���Bt�P��P8}���j-�:��E����Sjdf��Ϫۆ)˸f\�'��:��Ֆ���i���l�ĸ�'Z�8~�b�b��)S�
�Ӷ�N�H�,|�.������I�nkoĒ�o<�����\�Z��w��~cv��U6����\{)�_j������ͯ�xn�@��Ft���F�.*@փ�Ocn�|���%�,��P�xa#.4��$��9|�"�]���jz��X9H�Ț�VR^y?dj
�c�׻�BA��
�6{�}-t�*5���s�	�[��M�~cvq5ږ���c��Xs��t�Dx�v�N�Ǟ�?x��c#q�NpH�6���zl��c:9�C͓�γD�$7f;�6��"�V�c��i�-ń9�6[�3jؖw0�d�W�Q��N%|��_���O����`K��ax�n��ؐ���e��h�*��g�
f�5�Z��!�����������Iḽ�V��6%[�����e��3_O��c�k;�+�P�@߈ �����]S[�R�+����w��=�)%���fd�T7�SK��/Abpx�
�kXk�Gf��5�/(�х>+��6��م�3�T���,tD�R��Mm���h:M�N�;Q2�m���:�e����%���Z�{���x� &[���y�B���R��EE:�l���+t{%ȥ<S���|��6�L*����w�6ZO��W&&���&N��a�����3���a-u3�e��*����bE���§����U�*׻�E�/(9�#h�8���z���W�묢���XŤ/$-���H0%5h��o�s�$�"���j�>�zGY�ʋh��/mYp�)�
��}2�+����`��l�AVc�����>�z�w�����0���=�b��t��LG��6�6��u�=�Xij�
�+z���c�ۆ�[whB��<�]�ʼ`T�Z�����4<|\�Sb�YT4�=* M�� 
��*�=8����|�4?�T�õ�/�A�J)��@�e�b�X!`5��`j�w�(���6z++�ٲ���()뻇��͔4M��+�A>Ѫ���������Z�g�<���>��o���|�?�B��r�����Q�:Ɓ�8�#d�f5;)Cg��ҮI�P�����{;�r���\�:P��l�ҵ��}��2D�3^����#�
�Vx����<���M��5%����lrYu��ǾF��rx�v҃t�Z;P�M��J���bڃϫw!K�P)�m#BGr$�,1=�M��WC�Ҥ6���n�FF��(%��)jp�i~����]�����c3���'��K4�fL���1l'���_��[��mK��?Z�T�KN��2�)S�Ġ~T��oU��uZ#�i8a��w�:E%!�I�ԴǛ�����(OG�6��f�y_ɏJd��P�j���j���L&a�s�z�(�9�k--a>����JP�xc�:�������n�h�Dĭ(w9�I@�,��*#�_3���ͦ�\����
�Y믭C��2�}�����F�ꌆFX�l��eeC�=j�j��>�I��}�n��̟�v3`{�z��Jʛ����=}���sQW�^1�S�����
���u�ѨAkHp��N�H�)Zڵ.-�M���xQb'^��C����Ү�l�J,%k���4�]�(���a6ii��B��^p�Tӽ�t����ף2�}:��l�U�n}�g�	�5�d����M6�*�|�Q�ǶNQR:��pˇ��A�V�t��5�R�B�r*���ГШ}�e��d��m��q�j�ۤ�����k~ٗѸ��?�1��R�	�	�v&+>=J4���q&�dG|}9xș=���o�K��c�@�u�����ѯ�HD�O���m�E�!���'�N��o.),��)ݻM{,Us�!HWG;���	̄O6h1#��������*fM���nN|l�x���w�XgM�
VqinC\�Qr�S�I)�!4X,�� e�gRr�x��n(R����=e7k^�ڝ�:#�f����E��zX��p$6���3�b۰r)�m����Vhх����h�N�����U����-�4m��j*>ͣ�{��A��j岰���?'�x���}��hx�Q�s��w�R[�q����K���d�p�?�E@;U�>�	�~��Bٔ�K�r�SD��?
��2'"��R]R�g��
���np��X���g�sıc:���2~�w��h�3)2�q��F���x��x����ۖ�w#�7��3K�*��L�����t�o�Z�����r���Vlo�:M$�x?hE�p��1;E�G
���U�־wO���㬗ͪ4˗�-O��*���3+\�0GW&U��xo��<�m����V��~S���x�Ksӑ��+��p�q��� Q1�rJ�m���ԑo@,�R�Y\f``�]�,X�?���#��
�m���-
h3�s|l���/���@	�6��;WjM�q�B"��r��9Z5ݭiY*x�i̅�{BSθM���OE�z���	{�=�A�	zs�m����b�~0��-��:!r&ɬ"�um���w�^b���X�x�9�&[�u�za>�~EƏ}]\���$�3��٘��;�#��t����r��N��~E��d�����1�K�0}%��iBG���MC�U����˱�~�,�q��|C<��2Qk.���� h��/ֻ�q�$ڼJ�3ʋH���t��S�red��쪸ujd��8׭��eg�I�l�����:�K6��Փ��k��>Ƥ�����m�T@c��y�֩�MMX�K��/�y�B�:����5]��&g�w�����mq��N�G6^����'%T���{9�3볨U��3�%hg��XF�q�/�Ƌ���m�����e$��%�y(4� 񯋪N&�%�)��줮g����۶���kn2UvV������u�۝�?��@��3��ڂ��P7N�{��d������kfw�u���N���S��~ �N�C�E�'�>����>����9��T���
.�2�i ���C�М9�b�@3}ȏ�"]�5vR�~���IW
~5�KX�0(�>k�#*4�����J�Y4�,�b�m�99y��1b�
�^����?�R�Q̇]	�F�/�ΘWR*�V�������������Ju�P�y]��aL���?�ڙȋp'��B�u򢴣����淨�����*<��ֆ5"?���ύ�a�6�
�D���uR�U�Ѯ���3�ip�*�$��㲙�u�} y��5;��̓��n�/<
�Z7�ix%���%�},Y�9��,���M|��� �:�昸5m���O������T�ml�y��S�&�l�c��J�=�<��K��}�xh�t[�E����2������Ql�37_�u��U�.JgEw�����E��.��Q�Xjc@�Hi����\���w���p;u�y���Ѷ*;�2Kye��(b�`���m��,��A&�b�V��A�h\$X���Ҫ(���]��]���5��:�LZ��#N��X�K�[[���6�v{��Y1Q�unl(F��ru���������)����� ��,m �/f�LN1�ʹ���4ͮ�)_8Ь�H�W̚�߆��v�t�6�\+��fդ)�k�Jo��!�Kb��9��9�I��M�j���)	�,O��E4m����|��R@�_�"ƶ���g<�O�v��/��y ��κ���D�q�ų[i�U���f;F-��*!�>{&0�ڨ��ʗ(<Ŝ~�EB>�؟c�$j兒�h�m/r�}$���w��N�j��{/���NE��I�j����佩j�������vA4`��w�[�(J��RI��X���wL�ƻ�R{��KQ��69;z�Z%�Y+��#�C2�r][~D�0���?�϶�o�s$(y���P)�i/�T�ݏ&��r�{��"�xG�S��c�b��������jT��#�;
'6�ͫŞ�o��n�(��T�t���KG�1O�R����!Yq�~z=�x6� �{�����5��G�8)A�x�)4�u(}���)��\W�
c:�2�@2�f���+�C��!^bG������w	���s�%BZrh!K��Q�!����{��s|�t��P�{�X6�FaN#�m^Dn�Ŧ��Ǧ�!�Щ& ��[���.E�xa�d�~��D��U�����u��&�r���v7���:��ڿъ'���%n��L��xdF�0�m5��Q���k>�˲��_���z���9����ڨ��]=K�Z^��+���O�h��}v�3y����d���_��!`�(eDf�a�y���k�p{�R嘱k�6���<"�D�{�����əs9��B]X��p����O�l���l��*�A���T�Z��of�q�vH�����g��,GtA��W<��?�N��911�����MXx�a�����^�P�i��]�k0��B�ޒK�*{oR�S-�ے��JQn�	}Urh]���*Q1�b���LU��2a)z��u�s0f�����k��1�K}EN-�������&tX�m�_�l��^65��G�OFA�	-� ��*� ��Xa��-�8U>��� ��2TV��WD��kQj>�D_鷞�%';��{�6f�@�������! ��ݢ�
7��~�;�9�%{5�yQX��ً�'ى�����&S׾>�4�CSw7��06c�Sx�����/H���Vf2�G�e�Th���L���[7\�?���k��C��pٛ��#PG �H�?^Y�A�FX�t[�M�:𳌋O1W ��?��%��k�'̛����D�8i�0"��#��xN0_$ߝ)Ҟ�y���n��|y��.H7,M�ïΩ��O��*��ϴ;���lh<�C��1l��i'��!�z7�tԕ�ɯ���y�nurT�Ӧ�x�����9��n��_rº������]T.������vuؽ�:�Ծ3���D��/ɒ��@z5�� ��&�S�`��
�K�n�m�'kB�ê�Yy�ƚ"W~����Roc�E�cܤ����Ld�����Y�H֏s���#�K�]��Q�|[����)� 雷��A<?��-�Z��}�v����u�7��a#��Q)�Z~e��g�~ V�s�4�A9�\~���6�5;R�Uq`3�6��2���[M�²w���F�`�nV�k~�$6܎W�j3�%�^�g�[�)F*s����M�O���d=���t0��.�^����d׋��W.4H�=�q��כ�tQ8Dma������/�VP�����z�ΈԠIUv��J�R���f�H�����oƺmu�{v�c�q�fh)wf�JpZj��$�(��%<x�R]��JL�|��<Δ$YVĺ���Ӹ���>���7����3���b�C<��`��A)���m~��Ł�Ɛ ��t�Ǥ]��vV��l[^dp�$���1�2�`�l���d���V0?_�������\�����G���L��`L�X��J\ߎ�,�ir���T��y	�Y� �\'���y�w�qU�WyG#�pr�Y�H=�Ev'��&x�}��\�o.�V��gT{�"/П b@6�s�]�ʸ�v9����v�q����[�>��s��+#5�w��	˓�rzm�)eL�'��R"^N�~�LPK��W�LGANɘ<�X~S+�B�6R��t���i�-��@��z��\�?V8�:P^�{�I#��ׂ�b��G{��w�@���mk��i�5���q�����/�6[�ko�h:c�"LZ�s�(����tr�J5��P.����O����-�n����1{zn���m&�%�X���6��vP�����v�	�[4z5K��L���j�qѰ\_qW���S��Z/Mˏ.��kh;x�쉢�5��M�|Y(�C7н������4�Nٰj%�R*�\�j�ꨡ����#Q��Ie�]wF*�
nf���\���(�[o�!��kڦ"�3�Kl�k�۶��Zq-q��N�q���x�2!ĵVeC�a���|Gd�#E�s�?�����g�h�C����rp{�B���z�*h3t8\�+�ߞȈQ���P�h}L�x��⏈������q^4���.�s@Dv�P+�
��<A�|UM���4=*�� ��|D.&�,9���t�����f���������k�ˉlI��bS1�g��E�/�����#A��d�4�(�ea�BVք P.���u�;��ȴE6@\���^9e~�A��T
ؓ��y��2]^��Yg_��w���	~4�T�x�2B;o�D����E���;���S���_~(k��@���JJ=~d��""%m���۲ćxw�*���A	��GH�+��kǁ��qV�&qJ&y�h�ZhV[�i�!���
�c���F���\q��ɦ�	D�1�z�!��K�?e����Vmbr���s�d�
�FG�>�9���{�.�y.
��Y�R�"A�R'��͓_�Ž,vb7�}�RE)��
/�X۱����D}�h*�_�ȓ��kK�F��m���[P�Ӊzw/���豯1ޭ�ݹs��ձ�X][X�9I��߿�k��$���7ND��k^��i���b��ɹu��/3��Ԣ�\3�j�Q٪��a4z�����[~o�#8��߹�&�9��ShV��y�eu�$�h�)�L����$�Z_N����xu_u�.&�}��s���,}�%1	����cj��$�
�g�3�.�D�w�m{�f�:˗i�,$����e
'���L s�WB�V�2�AXȭ#�����}KЀF��:�.�E�N*������sKn絮�eɌo����\D�M�L�u���.Rq��C<{����7%���&y9���^�7��l.�_O& (2���=fo���ߪ����ʏ���ְ�C�^Z==ɩ�b+_�o����wX���{��%�V"�p=�Ӎ:�j��ݶ�*�b��]{SW�.{@~��њ<@��\��.+�g���<^�$H�~p�Uaධ��N�cq�ԻՂŔ ̕�-����l������bS�Z����.f�.�t���7���$c�C43�uw����t t�x��4C����D/%�b?-`Q���Wj��9��r�{^m�����m����6{��|�Nm�^9K�Rt�ˏF[ t�\�FsB�RĚ�#&/"��������N��F�j&xz��~c�O������U����Q�tr�]1�i�?OĮ芏��&����-��N�v;���l�\��z�#,"���">�{�u�o,$°��0���ő��S�﹍�11y�vH��N@ WUi"9Ú�/��pWR�>Z��;���~ʎ$�s��-�Y��J!�q6dE�;���8<��}P2)['�6���Lά��N��v�����s8.U?�׻zo|�23�W�W���{�1	E��\�G��cl�>�]��z���`8���no��%)���C�Ӑ�~�zo�Ѵ*o~��p}���+U����_�k"Hu5�?3r�66-N��H�J���=��Q�=�!�_�~v���"*�|Č(xIHY�ї�Т��\8q��y�ܹ9��OƉ����5Q�~�'G�@.j�-�*$��Q�?�q���z�/,��L�&2���̌��ʣIn�c+���wt��3N�W�e�|8�ͬ-�Ӂ�ߨD�>kS9�ߠ���hg�Y���Y8�;ʝ�(�BK���G�i.��?��{��d��^�f44��U!��i%������"�Y>��4�Gj��ʒ�|eQ�1[�����J�o}Y�J�q	޽m�&�|�f��y�R7��L{̽ךV2M6n�I>���a��Su�m�eJ1����?{�u31J���_���|�͹��Z��z=���aI'�@��p��աsMa	D�e���,���X�׷C��jު�~kܾ�G>mV��7�����3�L�z�!ogd�x�@��qyL]q���58��v��׀g�j��6����<<
4�v.-Q�!*2.����z7xJ7����M �॒����� ~���{��#Ϩ�+7,��9>~}��C��`��� %V�`z�;��������	�F�M�@p�<��������-Xp�w	���5�{����s�}�o06�ꪚUs�^�W,s���д=�L���wה��h�f�c�����{+��i�"�5�,�3���\��I��y�Nv�iD�09f}������sH�	{�F	즶�ܱU��c��2�t���S|΅�ҏ�|��w�(�fb`��{��0�~��P�v\?GK��cZS�>g��;>y��K��O������A�+J��>*vGA�J�������V��k���[0��
���ҢΌ,�����!���������:L ,�X+-���3�\9j���m�(����wu�Qb��:�Q�K�5�V��~/B`�tC��5���y^�CV�ls����Vr���Z}e��l�{�7���5�[\�cAp41�K���ۊ��kҟ� ��BS������g/��3�#���U~vd�?�����̋� ���M�/�?��7y���k�͆�g�����)}�	��!� ��װ8B��������X��,Ѱu)7߾byȺ\�@�m��,�f�J��sjk�6�L��_㈈�7?��@��T���f�;�$ +O:HE��+v��H]��Tu��W�iN&�-p�P�7%�'K�4�n�Ǯ������?�pɳD�~� �;�5�N$��Z�t8ﳮU.-N���0~�Gi���;����\��05S�=E������sj0MΫ�ß?�|�
j+�V\�ˎ�b��ₚ�HX��a���܌��&4�`�=N��L��m�i���i<N���ڪqm�*K���A�~�o��]�l�4B9�{(C��������B�,`�ҲE}?������Ĉ���#8ϱɻ�|��y��1�s\x�:^:bJIz�ʷ����~��աm�޼J�n�Ge���f��ǵ�^��"/(��n2�m�\�ƕSP�Tx��c�Ֆ+�9��NA��lB��'2w��{��C���F'�j��c����b���\�5�֒��X�K����[M��M}"5L<Lw�eR�)�޼F���^�L�B7��Ol8��W:�Mzŕ�B���V6�k�&%<3*c��\�%`�d9g�y�>訷��RYa!��n[k��&�j׉���ݢm�.�6f 
^�����B�=��4�&�R����D���fF��$��]�Z�x������uWE���ۆ�K���c���t��[���`sY;�ڽ�����Ѫ��_���M;���>��?�>��WMF���>ސ5M9zk�.��?�yz��^KT`�+��0]�/�q'y�}.*����:��,��i^;����
�s�������9�ez��ǔ�n4n$$R�A	x�w7��<?���kTap��2�}d�"!��&�0�VEN��������i�d��>f��L�ghYY�9rO7���{�*	U 	]�\D"8t��.��ci���&�YG��Ύe�$P������w�,�|�b�T5������]E���֕����@�*
*F9��:�5�?W��]��0��dr5���G"q�A�]����9���*-��P�ni�^���}F���\#��&�q[�Lr�2S��}p)�y�E���|�Vo��a�RV|*��*0��M��¤���5x�y]�󭉭��·C� �f���(�g����Hzv��S�8���bC>B�v+ʹ���[�I��E��R<���@��ݭ�]լ��w�a�����xߠ,�<�a��8�3��3U2g	��V���������x堵���:h'kFB¼+ʨ�����
�[��N,���ޥWGT��\8��*���auz���O�:��D�0�K^BХ(�[;>!̍IC�;���tx��խ=)(<b�Ń5v��3�@��}�u���n��K��U�4c[�5rNӦ�L�3��Ⲃ:l����a4u�ۨc�FX}�U<��C�u':�xu�{��$���k~%�4 �;��@}�ʆ/��	T��v�:fl>(-}�D���|��y�BXl��K� ]���~�R�M�<>�.;��Z�U��[	 �br�NEF�>C!�P�������)}���r��C�3��T��1)^��T�n��-�t��Ʃ�X�E��Ï��J\`��fp���7c����$���d�H�|��0��
tm�+���T�$�vqD2�Z*���fD8&D����Vݩo+̲'��1�$�X���	����g�M�ǻھ3s4��Ù�&]8�a -�Y���\��#�"�.�j�h��'ٶ�M��oi����ή���^AOm��-��'�����'���������g5`�O�tE�ޫ�XPн�K��!����ϼ?���M�»�K�N�%k>��]����[_|D��?��HD8ؠ�+�Ҹ�D A��&��)�S<�?<ZX�H�E�"�T�m{^��S�[���K�qmݶ�D������&�o�fj���7�N��s�:S�9�	�}�d�4=�r�:ij���5;� |�%�����Ƞz����j��d�Wq��$� �a��]_���\zg���`O����%�	�c8����N?F���$kT,m�B�s{⮜����n�]#(,�bΨ{C�{i��Hp��c��F-J�BUm���Ad���p�,+�gz��۲��f�ju��XlP�Y,��[D��1��f>�8��
�_J�nS�cc��3�V��hq����;��}$�TS��8��������@�l<���ېL� ";�o�,�� <J66�3 9� �ǻ�p}��O[�E���R����#�8H݅���c���!yM�ڣ��ބ/N��ҁ�ٚ��b{P���2RRFYA�¯G�8JRg�]3�;b�b��HS?e���5�h�m��IO޸c��ۮs&��uaW����l�S7'�XS�����;]7�m5�[��g~�ccGs��;�Q\�ug�e��Y��	6Z����n��4Z��
A��I�6σ��hѿ���ߟZ���=����>��让,��}��WФ#`bJ{+����,����HL-l�;�1aݫ,$ԑ��5|�*�e�צ�U�lMX��� �R\ɩ�]\e5HC��_�*j�+���Q�}k�+}�7#8��d>jJ�q�?Uӧ`�:ɷ<	�s��1t�`[���|�qyp���'�@���M�|Z�ek����!al���2���;F��x�AW$��l�E�t�թ�����K�'BN�z��O	 �+Ub�Ԥ��a������#)A(!K�أkĖ֘�N�7(>�D���g۳��BS[+`�n�H�4�dd �U&2��6���@�ԗ��x�åL���ȬC�OD_9��8[(J�j�1�а��Ŭ��_W�-��B	���i?&m�>/��4k?�1CL�Qj��A�ۧa���Q�#{=]����jy�G彘#O ֓�6Q�|ڃ ��Zj�|T�(HU�)z�)�x!jg�#*���[cc���c]�:B����.h�3� n�܈�H�`yZ�������غ��N����^�mC�Hi�����n�;�\WՖ�� ���T�Oш'�-�k����gg�U�K�ZՑ����܉go�S��k��2�����@��hX�
���4s�"A�H����R �'Ezu]�P��]V�4а�t��5L'vUJr�� ���?�)�G���UQ��X���B܊G6�S"�A���v`�B�=2��&����6����Y�b���>�zm�>�VK<��8t�$ xL���DqyIG�[>��*"���[��\=3�s]�#����!
���ښ^Cf���J��0�mU��q*����ك���>a��s�ш�I+�V§ ���(���L�GgG�5 irT}։�j|A���JW}@?Y�'㎬��X�\�-����_��>,3�n{�p�>M��SC{����R�	����GW���G.H�;?)��H`W�AC���'��{c::z��R�l�>��Բ�����6*O����l��A�O���Y<E�9�Rr�2����s��ɓU�OJlt��=���lvo�Fyyo� ~e:͋76�Elq���Y��t�,B@'�L�GX�A����ww���Us�T���t/��[�Oi���Уl�M����%,W�@����^���d1��kz�#��ǯ�k#!��rN�@/�>Ѻ�Ң�����sk|��7�rS��=�0�y������/7P����#�!"q�Җ��C����[[���|�'a�̮̭���@��k��w��<���|OP���@��U�������jچ�n--�t	�V�U��+;ې՟�0z���A�Ѹt�ܼ��R���ު,NmG;�Ӂ�1�����j/�OcT*gR6�0�HY�a�����}�u�x��2���-'.Z�f
/����Y�8smu�g,Q����?��'+F=���@��!A+ȳ
):M������[�����I����	�*���U�5K��6�Jut�!��F��p��M�k:���"�45ß����5��;���脃� wE/e�0�>�Fʅ�O��m�_W��&��U���B(-�l*"'�`I��f�G��Sa��!ԶT~�gHϡ�di��84��sNlG���0	,�<N��5O?��>��++��kQ�T��]9��}��.B8?�wKTL�lt��\u�-�}��M�����u��Y��JAv�4������B[�큽(�\�[�Q�EE��R��[��}l7BO+yV�OC��"6�ϯ��U/��"�~�����%�3FB/'�o�%c3O��wR�*Sd��)��><5�T˵-��&g����������F�y����=�7�(Df�d�t�L���{���
U�͉RRVw������C�ĥ߈.ɽ\k4X���/�X���Q(����"d`��ݩ,��PRR7۞�KIMS�F�rJ�$G�ڶq�~��9e�LU
SV�M��o�FoW�ł������_��������?m��G�=��e�R��Z�w_&����>��ʤ���J���^.�����os�-��&V����2�m����4A�i�i �$�.7�gש  |��\A�5wȊ�!m��q������p��M��V9� r�bKx�I��~t�sp�ф9H{���lֹ1{�S)�d�� �.�z,=OT�	�HN��(�����g������~����{O�?�rs���uxr�;M�Y�����5a�rc5�%Zh;�h��v	����6���[��a`�Բ�w��1�D�������&����l��{4�6ψ�cbv����GX����p�OU�a֓1�շ�%уV۾��aŐ"XFQ��ۍ���-]��X��4is0XJ$���&I��K�j&]�����~���h��Gа����n���\l��R�OpWR���iCܡ��OeM��Bd��Z�Ñ�bj&F����P�0jqҮ��r��#6��,x���Κ8� �I ��1fE��������Xc��	���"�5���5L�خ�K�k�%޴�cL\��8 �|�����>�@�;� �Ya4��J����J|VϏo���=��$��(,�Y&�M��ς�@�/���>�θ�l�$�؈H�o�V))�����.7�M��h�"���6-H|�}������D~�����V�SN����G %:`��k��x�Q�zy��B22do�1�E(r�Tq�^B+�Tj�~Pv�m�� ��Ғ�f*�K`L�p�z�}�?�s����D��v)�'uI�����X�l ��G��I׶���N�d�́��#'hC����͔�u��P�T)X�>�g�x4Gfs'<�r��g�b0P���"pDO���}�?#D]{�hr�Q�{%������X��h�߈�H{5M�Ȣ��"���F���gK؋���t�C�(�n�ն]��+�kGV�ި�t�Wx׳���tU�nS��ocՒ��3�o�p[����9G�[�E&f�������́��G����y�{r��f� ��/��@�O�;X8tq���*��-��Fs_����~������6}B[��&e%.ra�����Ť; ����}l��٨Z!�:|��i�Ql�ޱ;>0�;���?��p�����^��g��gn\�n�DS�ͤ�H��]\8E���u"�df�j}hLs�4�����hkw7}y��Z�$#f����ގ5����x�aBl�)��\R����+ U�[/1 ��U2?�S@H�=��|�~���������y�����M��S����Ԋ���$�s������*��lqA��LH���Ԯ<aq���;�Rg~�,��e�-:v�cY�@�]U�G��+qEJ�x�_}�a�\���F}ߵTTb�暗�y&yŮI�K���!�:,�=�wSԽ���P�TON�>�����)��A��K�ۈ�����|�z�>ؚCe���9����'��H��"_d�3@49}}��j��g�Y+�`D"����|)%܆���P[nH�����s"DD0TJ$�C�����������x�'����oCC ���^�l�����|��>$�,����]1�{�X`�����q'x�ʖ�%<ڝ�b��/\�����]N�r�ַ�@��2�I��&l�z��ֵ��v��vh��Vtagb���{X��uƷ���X�-s���ygR��5���:˄N[	
�;�e� E����1a��1�GP$MI!����"5�H��Ӏo>�w��ۋpwV+h"9�	,Q��-������:�")��1�W؟��qc��@��H� �Ny�+��\�K�m�Ѕ�2 �"RJe�(*ﲰ��_�X���
�K軳��	]K6A��Y�7�Z��R�0 �]GN5<xKg]�o$�nL�F�J���m����oP���e.1T����~��j�,-�
���}u��!��4	�f�&����Ǿh�"��xl��6�N\7I1��(�]����^����`b~>Y���-4��0����b~��1�\o��3ޔM��&���ɤ����M���JZ���l�a�����}A���I87��9)��C�.�{��s�5����jA~�
���)�|�Qkx�:Pk�DH�b�i���=T2S��#���H����]����9�	������_��o4 �N�rԡ}0&�uy3+z��^b ���e�),hYG��7���$�zI��*��8�ґ�A�Z=�րp��>#x$�U���tb�����z�w�ޏ�λo%��/;S���ZX��C160�$LH *萳��r��C�%*&ez�
7>�FÔ�)9hav�W��������g?��?�˸��.�������eB��e��J�ZW�n;�����M�[kW��!P��l9-ו�ph�K�f�T��h����%�t!�k�|!@���у�.���232��|鎭������Y�BV��-��f)��O�A�=ǅ��ߒ�:���Y�U��;y��~ lԀ-y��H�4�Ofj�a 9����kjޮ�c���JL(c�����ydbd��P�5%�gϛ⪙���5���S�jǐ�?��P}2���¨-������"��s�`���-`{Y#{�t�E��6$L� �8}�Z/�؝ �FiII}31��̾�!i$��k���ǈw_���Έ��oQ�B�8Ɍ�!|�~����G}$>fʝV��dMf֩\�#��B��̏p� 5q�a|���J{G�5[�;�B{p��"��Sf(���{���}�4!����9Y���LE@@��^'AY��	�C��3�z�f8�K��V|��yQO�(�z�u-��� ��+ZZv_e.(B?���V�����Cg�t������#�x_���f��:U�f���F�4ڣ��J4���q�n^3�n�����*]���1�����@q����Zmm�[c�{^�V�1��j}�{c�r߰.�}4�8���k
�EYN�I M+g���a���i�da��oB�(��T������`4o���r�����8�ڤ.|8Q]{�-����+F��j����^�Gl�X�f>����h�� 8t<f&c!�V��ӓ���dE���F!��!;�J�XY�t3A���X���)&po�h��8�9�Ox���+,�@�ܩ��㸷���$'����kN7��kh�P�)�_��@��K�A�9ܴǟ�pUl	�I���`�,N�a�܍"�IY[=���qi@�G�:�N/�?iԴ��P]Lm�W��U�%�{ݟ��?T��ѩ%`���5�>�b�8�[o"���`H^����-��^�z����b݋���~�i΋���Y �ΗhU{x��!BF�F?��b¸_	��.N�
Z���v����MW��9Xm��O����u�H� ����s):�����(���^����y�:�ti8]���:8'Y�\[�
�¥BxE��n*�2��/Q�5�XZ�]$�AlG8��u��t������L��25M�A[P�}���ۍ��?4�#C0� m���v�1���,8��/�������_B�j\��,D��2�i�PH\��p_u��Lö����"�QE22���s���.=�'#��ɮM�q����Gv�+;�'Zf6��ֳ��ut�}��B��|e8�:���űNWD-�'�䳺H����:�S�b��1b�B��H["�6;z޺ ���uh/@9Y�a�l�#�g��^U/�F��7��[�rlУ|�����Ƌ��m�
�|�RC��k��:��Ms����|�&�����N�x�8�1K������?{r;�i�^��=�y�Q��S-9�W$T�|c�:׆�!0�W��9�V��!���xmKG�Ah@�-�LElA��?W��8��b�� 8-��v���8䇿��|�Rh���&����QS�EAw��t��"ц}���#��)rmJ��m&�h\������W/�0=�����N��ML�O�P�H$k�H��Z��&ī��8�l���*}�����&�+Q;�
� C��?�7��ןLe��7'������s]���~2|�QT�h`��h8�OKK�bK�n�� I�@���������K�!V�f�u^������~I�.�{�q�NA-��j_]E�7�`ωї.�&O#$!
'jId��'�t�-����;<�w����s"��>��&#��������q	3�`�dl�ɶ0M`L��>)7wD�W�����z�O�涎�3�n���-6�N(�y˺:���<?�3�|y��t�Tמ�,ڃA�Q��>��+cu3~3&�zP#�	}��|��m��EC��,��l\}Q�R�ס+yû��LOY=h���eq�>=���������I#nz|��l�cib�N�����������**�\g��"�$��������F��@j�_t���,Hn�'��޶r�gmϾt�<�\�}��pS9�&�gVx��B'&��oWm�V8����NAǴ���[�㚅>�9����5^܇�mo/N�>�M�_D|����ս �('fF)��RgY�>��Q��>o�zz�j���W���{�~:��'x0~��)�3(r��7GΧj��W5���
AjW{n�$C�+E}#���LF�`�,��%�����c��.%���J|͕���c����J�ЗI�j�
����O��UB̝��~7B����Z�J9�ׅj�o���"?IZ�qO����y`��i����ٳ�/��), �S���c��=�p�_�>��,���z�Q�,z���U�evLX��޼�v�Np�f��ni~���U�qxr�ے䦄�Àѽ'C����ff���v�n'*���P��VZ�Y%q	L��.�G5������Bh�Z���?�M�^�*~� �D�?�+*t��-un�Q,�D����!y�d���.���-������Ҋ�t��/�@���AN�r��,44(-�����Ǿ;�N	��M?&�*������"��S6#�r
�����ך,���f�����ܝ>����胡8��0�B����{����>�X�������������r]�~bCsV�cI�!����8��.���p���ݪO�}�`�C:�z;Yy{�#֬�"޿���v�,@~@��)�"�ZiՁ�Vpp�����|��Q0|�A�R��x�����(�����ϳ��nzã�B��P�v�F�y�^�i�-6�&n�V�N2��O���F �v���IP�,d�GDV��@����=J:�Y؜�Ce9��k�E�9�c��e�Y�I�Sڂ ���WM��)_kbN��HF���y��-�����+Ψ�P,f8���B�v=�4��GG�sؿe�/�$���Č�Yp�KK��T=�Z�$v{]��U��=�R��	3��6!�}wo4�#�;��U���Z�r!�ؗU��]��)�m|���;y`;:���$�̄Β���Ax���j~~C҄fj�N��
9y�8�QA{m��f�Վ�*������ ̓�@��e�ju0�!bԁ��B�K��(@�PR�l���
���� 	�~`7h�r֙�\�8r�5�L����1�!�e��,3���C���N�ِ�֦=�{AG��9�ƞ����!05�(�"SE5"�K7x���֘���ƈ�߿���"��i;�	�g�P��/Z��R�?�뜽ؔ�MN�D"0�� \�Pm��1!�;�
�3�M��g�7<�9���xL�MǷK9۞�M��v�����-���R�wu J�Q$��OWE�ݲ%Q9���|�>K�Z�ҏ���0i=V���~{"�O7o��sV6&���i���֎�e��V�?�p�`ԝ������	����w�8�"�h�� �ݼR:O�w�.��z�;�OF���ہ=�j�P��F�`r4�^2f�f��¢��&]��p�a�YJj��r�91�
���ϼ���b���u�2jj��m��t=;?�mm�V#HD�ڷ 6�x��{a� �w{���r������F�����7�\x�M�ɫy)iH���w:IJ~���L�^�I[�K$�^�=�0�w�{�		f�{���
����Q]��>��F����=ek*|J��;by���A�	v��Z� ��zr{��'��1XXC�&+�zrڄa+����`a�݇��,U!(Mף���{1�^3!�f��i<a�?K��5W�xo�1m�\M.��0����S����%��6�Cs1�8��}���-@l��>��B����#�qJc�%���e���xI����pɴ�m�uI�Jx=���Q�`L��rH7�C�ֺDb��g�k�
��;M�C�~t����պ�#�[�Ok�K��"�A��?�Z�|A�eLcx����e�-8a__�u{�_�C��S�pfʘ�G�w���:|����6tl�@�>`J��W^ݖW�|�����tKk�����Jnu^?�#�N��џ=�|�
�����U����GH`w�e':!�W{�3n���H��-��B����cc硗��Ȥd��Q�HAK_�,s�4%����v�|p���膮���q'�����3ʦQoT5FX����Z]�(2�Bx�biő[1���Ia�xt)lY:�ߞ(����s)8�i��M�?��w
Z�ÆZִ���+��59�?�������d�W{�4������G�&��>f)P>�ᯡv�O��46Dn���E�+�s����	!l&܀�
a�"�v�0�J܋�G�J��\����:��>3p7�柬�H�İB��ؓH[�����y����&�{/�ml� �'���_ߔ�Z�D���d;������V�Kz�-��8��v�N���[���\��M�M��u+E����ˮ��T,�?ѻƶ�ç>�˞>�M�b���IL�\���O~��q;��5C1��,��f2a�>�Ǫ�~�|���SE�L�?M�c����˝/�js�Fs��˚|X��]a]�"�ow��vqG�-�o���Aej_{�tsp�\�U�V��OwD�����:2��['�8��S�|b�O�W,�P���;fZ�Si�?&�L`�+�so�~,.�oz*7�AVL+#p}��e�J����7aXd�Aj��rh2E�\��2���.ݷ�ytM7�0dn�2��t[8�7��� A �7�Y94�a�O�"��n3// �0�3z���f���2��&F������b��ݻ�S�F'p��!���>{]�h-��Z�E}����ɺR:OY���Bqj�4�]GL��sN��LP�4�/��vS6.u�{r�g�Pu��C����/�w���noK�T�9��;�T�ʎ�)-���6�4oWv��=N����`����L���5���W�0?�@;�Z<ƶpۼN��*E�n��j�"e�Fʙ,!Lx�l�oƃ����ٌ���V:��\c�7��%�r��ԯ��
"s�ֻ�e�B�᮪�ᤒ��h8?��#4����w�Tp�v�ړUm*l�g�H**�<+;T�y�$Y�Q��uNo[%��0nt��o���e�n"�Z<�++Z�����:]{�Wan���#���\���P��E�|r%�=��'�~�qT��_�,L(�������(�vq8F�����Ͳ �V�W0Ҍ#KMM��Q������E���L�n�Y�:?�����r}��W�V�-L}�aq)w��!9���N��|>�籌ѝݏ���z�e�u���25���bbVe�?]eS��q���DN@�[�/��x����7È]t�r���s I`,����16���|z�0�	�9
ƫ��k�V\�������0Ll6Nm
�T$^��v�U�Ub@i) ߭2pZ�E�HH`ZuF{!��<D[Mă�����OR�V�)W����WT�U?�<z���
�#E��ӴffJ��&����A���ۚ2ߺ�O�l{7���ڨL��i;�Y�!7�����l�{��->�i�J`�e��)�͇JRADDl8�\[�jk���� �	
ƹ*@z��"�-�x��HX(��>�rN�wQT�^�
������)-Q����dyώ]��ӳa�Ѕ�|�2 z�nba�eJ�%G�6;��zކ�/FB�ܭ}֖KA�nPg**#��z�1��p��P����P}�oo�Gޯ���d�t�R��
�й3�g�̖W̙����ƿ�SV!P����o�VZ@E���ۋK�&e�±��OF�eR���hS����?Md'):�v��4Q��ɔ���U���ѠlrGa+rJ�̺.%�P�1.�L�l�2�:	��T��+(��x�	���v9{���6��ü��k?߸m(�[}�C�*���1��j�C�4�d�����|w_R|����D*�h�I�m�hO%1ѣ�(�͇;V*�8�gp"�ҁX�7��D�--ïmO>>
�21�2�A\��Ԇ]u���J��?u�2`�]r ��^���"��RBK��_in���C;�@��*�9��L�O�		���2�俖5?9�0j�����g��)�W7�,-�v�I1a��k�֬��,(�>�p�޽��C�V�V�isSH��,b}ɤ�YC�7 ��Isaj�G�ٵ����0)�Ej�𗒇��ǂ��^�L|%�,G��]���[�,;�3�Γ��t�G�-eō��hڶ��j��w8"�4K'&"�0���߳�J�}�{�h���thҭ�M[h����4������.J&o��u5K�p������^�<�Pe�`Z��t3�.Fi�Ek���o��hi���
��Y�>|PPT�����(X�Bp }��[(��^�ί{]su�Q��������"��.)IsK��G`��̒�qE���*+%<�2�;IB1�K�\���7�'զ�
 1C��5Ks}��us� r�r����NI̦�NI�R58��A�Yt�Z��������יضh�Ϋ.L�Ah7ߥmr��H%�+�]E�S� 4R���^Ӊ�vj��+z9,ٓ��'K�����*�=l��N���E\<Р^���l��?�p�|�5\�@j�:ɺ��tD2�U2y��F8x�c���e��A44^wZ���g�";}�ejX5�ynަr4q��4��@�o؉����l�,4�"�<�X�1U���8��D��dEoՀ��K�X�3�cY�|��L����A�]hP+����k<�G/��K������^/NQ_�X�c�5�y�����>�`�Kޝ�}��(E���nh"^Q�)�.�ú$�!u�KV-�	����ݗ0��nk�xWy:�x��`?Rt*���~���r4$�]�c������ܶ۳T����.�B�ͨBkS�&:�/));���#&�T�9q)��ʼW����cє�O-�V���������i����2r�۞�ԗ��**�5�Y=� =K�є��E��H���Um��fV||>?��Hs۞N�`ݙT*��2xjWmf�zԱ�����ַ뱼O�R	8\)�)�0n��|,�-[�������5��(�Cӎ,��ٯ��[ @Ȥ�eܧS�i�[h��ˋiyΫ���ѡFFM�MFi镪>�[�?<����xw[!B ��t�[4��&��ͬ�FtJ���������h�7���q�ʖ18���s|*p ���s����b�!UąA.-��Y��i�+��Ï�-J`�&�+a�ZMϔmg�|=���L��N�ൕs�������!��ɝ�|�����֚W���rAd""�	z@pv�wm��	3�'�j�]��6�+@<n��)��by��zd4�EBW�����v?�>! �lZ9Zp���։�����~$�_�r)�Z�߉)`bg/�.-��bVP����fqR�ǀw&�˰B�Q(���|~9��s�����GƳ���t�$��"51Q���|8�7vA�/f�UR����vM��+��%q�C����O�2�j� �N���� ���L��,�Z;������Y ���Gw"KiJ r"� �UKl�3��k�-i�)�ڷ�o�����'�V�K���I����.F�弯J\m��~��?K�EN����9�V��¨@���T껮�wӷ4��y�
�HG��@�~�w���z�V���.��L*�:ї�d�]��~���Jª��3Sd����/uz��2�R.{v@7,̩�.ts_bj��gPFЋ��(���de�=Wb(�Z�̴��*d��=~�����/D}%����Z)_<�e����p��$_n��V�x�~�����B
�7�N��,������1��#1��%�s�����H8WY(V�0���w����쥨|�Q���l�$񊄬�/rp����������7:[YA��BI���� �=(��J
.>�pdD�چW\m��'J<l۳��~�7V����iMP$(�jKK�E���W�QR�ԩ���iġ�	��u!��2��_Ǎ�8�� �s~u[{��4hqj�	����ul���'s�vϡ�R�S���,-$�jG�5rJ��ѳ���o�ܭ�Ot��DE�/���ZJ���S�l@2�$�	o���<��7��>q�:���H� �4�DOK�K�r�NV�<n����9B��CU��1�u9�ǟHJA�� �q}t?�ç�3^<���ݒ�4��������<�W_ܯ��sM���*�����2� ����N!��/��b�1�����׊X�3����m&�Ɩa
�3�+�)�١Ӯ�������SzS��;j2<���E�~i���s&�E��PT�`]Q�`'�L�����XJ�_-,ʖG��Rɏߖ��ɇK�}8b�K�f@�(���Є����.Y���^`]?�u9�/����	^o���1�F�ӾRT+#�D��n�pL��h��g�Zi<�~�F���A�.'�k=�����v��]}��A^�&��g~�"i+9t�v��q�z&ŋ�:9�\ۻ�>������ay��K�y`9��0�-���d���뙼��f�99��ʼ��:#�� =%�iK֠,\j[�dd<�Y��*ڮ�I�sa��:&3���Q���T�!2i.��7y���IW�.W�y�������XZ�Cto�c����H�z��޳7�Ásۦ�X��k,]��&\����-:0�
�zO3+��h�i� >P�����e����K�o����ڧ$�Kf*�!j�E��e�E_������g� ּΟ�@�|;����Eg�k�Uc&����V'q���4p�M�:��+��ߣv��zW��\�B�\�
�S(˶�SP*h�M $���5!/�;�|r�[d:CC��l�3���W�%�b�� �}�����̝G=$ó�� �u�#3��|}A(a���p���#���.��1	/�t�e�}�}�G�ܹ͚T�6���.0L�!Lm���U3`��W� .��j����^s���;8��¹O�Lk�=�u<Q�z����>�]��aV���jy��	��4��=�O��f
՛�چ�~��M��J���H6J{U:�F$�����$F�H���
��G6c��L�� ���}��NZWΩ.r���RQ���:p��Ǯ��Nm�o�<�>nq)�Ғ-�k>G���w��Ɋj�d�=۾ڣծ�b���Q�Tp��7�>cھ�0[ay��J�VT�,yY���[�R㿽ȍ��׬��if5�R�r{;�ՕI��:�պp����9:�x�g���<������e����?r�%ŋ�H)�2k^���5��K(M����/煊"7��y�-�����!Y��]�浛����uhRG�b�Ӯ*�2P7٪�NI�����w�m�,i"�r�[��[7"��,�OZO��o?���٪�x�-�!�� �� H����tw�t))%ݭ�tw7H,��]o������fg�w�眻3��G�	�j�����J�(�ɱ��"&],,�0<�E*�~��������� &��)�L˵����gl�<�'6|t�w���Eb�=&�3<	�]
W�m ��1�%��O������1
~�5~x��mtH<�dz���}-z�.�f�?]\��՟������ک����q|&^�qT��V�mБ�LVT�)�quJ�L@�
$��B�"Zb�wȑ։�c�T��� =<�MϰX9������	K;�P'\�E�i���M]^YÇ=�EDd���#� ��}b�t�/�����a��V�+ٗ�-	��;��\N�Kj^�ly�&�GG��ʝw�rG����f�bM��g��'-���4NR��(�F[[k@�����e<l�\~�")���]�T�}�����٤�$_Ԁm(���g����J���Z|�U1}MW۲;�ە7����5����#h�#�PKJ�w���:N�f��T_�X�(�݂՘[����/���K�**o�]�e��BS��K���ZYY�(a�Z������_%��gX9�<l����c^^�*��̏�s��8�XF��8�Fv xg����r݉9��.}#QF'���ޫ�Mʹ2z�`Ä́��PF���?;Ĺ����8mŀ��p����	\f߆$k�4��~ǂmf#�w(�&Q�X�0�JCJ7-��a%IJ��ޠ͎|}M� �Ƹ�3$��5��z*O&SV��zp�%� �y��T����K��S�80�T��N��g�l��32b��)	8"�s������- ��5�h��4��뜅��f���f[�*"Rc�4�0C�nm�V�b�h^�ȣ�hy�^����]P�";IF�=��8���V�4ˏ�ζ��31�g���tzY�Q����&��c$8�ŅY��-_�Ѩ�EDGkkzhb�!�,���ۡ���i��#2IA0��nM|�f#	��hP�D�d>
CiF�D�%��;|�\�}���9_U�������T!�%aUe��t;�{u��S<0�
1X���/g�8J���\b�;I*�$��3��2%+�"JP&笞Uj�l�TYo��S����T�����^/� S�� �49)��2뮑���%H$���;�QCA�k���uX�V�7\԰�N*ϛ���;�A�V�ѲA�սV�i��m�&0��aMTaICF���4�w����W��;P�y���ʹu��)�B[R�?Q��N�!­�p��������ْ+���~��%l��ƕ����B� 	��E��6����Q���O���T'Һ1�^�p�`�m��r!�,y��A�p�bwI���#�??�-N�ѱ��N��u�W�fX~n1��X� �}9����%�����ҿ��E���v&^�����P�.KPܼ���'�d>�}]	���N��0�4���p�B���E�p��<t�0�������onn����mg[���Iﮘ�"���w?GAFqh�`�ٵލ������E���
��~I�8eԽ��)����d����%�E���=H2�u���pT�m~P�(����I�z�&���Z�v�V1:v�w�zS�a��,q��Ǐ�6�ۭ�����o��S�/w9H�9�ֶ��I^�$kꆚO�0MyeuJ?a�rD�fW?�,v�I��vĕT����� ��.�^��Tx����9!�r$a��tډ�Z}�`qЋ2G�}�`z������m�lh1���d��z4���fE�ٱgW�̱�d���F��_&��<��V�΀8	�F��j��E∁�l�d�9eu�Y�AW䤂��ܐn/n�1c�˪����C6��LN�GX�ǵ��ş�f���oPp���o=,J^��yx�0�3��`�a�!�[���|���K"��$����m�����X��GA6,l{�l^��r#E�ؖ��2��u�נ���٦��*�Vs�J� g���<�+f55�/��AQ](,��Ua�Q�Z�(�Bc�	��5@P�䢞ŧ��ad3pP�<@��h�	����!���d���W$ʜE=�O[c�R�Yi�����w�z��Q��51�~G��E�)3є�(�!��\�xm�&�d���M�;n�xV�p�`�PǀM��=��O]�F�E�M����p��c�}��z���C�'e����+O�J���3	g{���������`�,����l�+y{ KD�.�s-��]�y�k���q}�jhqLeǁ��H{E5�������� #�/�ҟ�WO�%�npr2ǣ�՜�H� ێ��*&s�{%e�����F6$���_��I$W3�E�^(f�=�}|FԹ�M�W�q�Ȯ��:�"K���N�����"�]uKl���8�*��F�Ă!��q��q��,�:����Π��=�Xj�ܚ�ڟ����F�{�7�%�g�[9j�M&���G+�������ې������
��{�Y�j��a����i;��ZJ%A0�ʀv6���s~��7z�N�*���?�NÆ}f�-����1p+��iǵ���f�R\D"�@��짬L�EۿS�`$�ue��6�* 5�G�=�`�����t�~�Ӷ���˘��L=�S�g(�W�2��}/O!#RA�!�V-g�_�q��o���Y�������� S�<��i���?L$cu�@��I� ��1�
77�?>�v:���}�sl��n�����a1�t��3�cˏ�6�*����#]�'�0�]�*��zY"�L�Í� E#���>[�4$o�0�m!+%�)�.UH���K�3�04��TF��������@� oX������-u�+(ɶ�Vs��Ųt�]��ڜ	�A�V:����N�-����Gב[���?@�։l�O�־�?�{����N�"�"�����x;��K���^lT��� ��.à�1]n:LP6ݩ�Z���0q�ᄰ}'�L/����AmU���]L�L�ݫ�Yj���04�rS(
�~�p����6й�_�D�P2�1\����=ƅr��,H����Q�I),¦�p���r
����j�$'��o�WC�o�;9�a^�Q^� ���N����j�(y{]�χ�22�i��Y���|+/�+۶E%���Zg8������w�q-�u���h�G_ʗ`�an@�l-V����:���}���$���c$_#�i�#]�?�h0���Y:�oV� 0�b�$�&�Qo��GFm�U����1K`���3I!��N���o����Eޯ�B�T�ǀ�<4������ݫ�j��B*����ɌGm�AP۵�z����P^Kp˵�H}���W-AO>��o��X��ò�o�h����"���A��f �r�S>vl-g����&���ň
���:��h�m�͛�<\���|ϗ�������-�݃�!1p~�S����־Y��c]ȟ��gf>�yc���~wY]���śW��kh�H�f�:�n����CQ�LT��������[�!�cK�G�F�D�։�����&@q�t�ς�Χ� �]�
H:�J�㯒��?��k��Z�����J��[�����Y�g�&MӤ5��Y(�-�8����_�`&ѩӒc�$$ba�̰�mo�v�/�M � ?��y
��]*%�;e�ioK�Y˥$Keyy�$h!B�G���#�z��KtGA?�/�UЎ�V �t����4i�o%*Ąo�g�'��89K&H�HO+X$OJ�Γ�J�Yt�@4�s�7)U�y���G1�ۄ��?�u�ml�	�~�������j��0 {��à���f�6��=��?,�z�To8�)�;l�C���zUy�UP;c+��w<�+�a�x�M���3<���#�Vǩ��4^6�G|��q���|̃)CH		�_q��B�e�*�X�����:�gw�E��'b�2m6�0��e��N��<a�~��G�?���[��Bu��^Sq��o���*S+�3�>n�l�V��jϫ�ȧ�����"�8N����ĸ~�6����+�������%�]Q}vӌ�5��DE[7xX$~jt�U0Mΰ��p���#x�\�g�����I*���?{���v[�Q��cVm�z����=bUd���ܨ4�k���b�_�Z��&%�,��)D,@������)-*�2f�����o��Pו�ʳHy_u��P�.����d�ĭĤ�
E�<f��[��[[IaE����`��o����xi�Z8�d�B�D�ze���O������G��5�����V�i�z�^nlul�{0[�
�07_ǖ�M�_��kk���rp̿-��L"o����� �G�����t��M�yl0n���>/K�g����1�H�"�{a�o��8]��>[^�k��sB8��[�n����A�1�MO�o�ۮE��V^�A�� ���-����fIؗ�l���5��Y!�܅m�z�$@�Da�\R����I?%��Dy�o_0!������uF뗩����]=�"u0�f�%��=�"�_FF�u��@m$l;�+�!�/b1��f{U��yKkJI�nm����,���K��;�ëQ>�6Fzkݎ�R��"�+���nf��Ʊ4
9��lA�fzz���`Rߡ��B�`FG�z�c�{m%cc&֭��g��no��xB�1����Q]��:�8��_:���:�"`�o��4�m6f犒��j�[A�*gY}��r�����̾���Jc�͂IEU�Dk�O=���P)�T�W�s���w��*�cg�?�	(.���q��U�� �����;F/�N���V�Bg�FwUNW"���@�(�]�4� =�:���꟔WV���m�,����i/�_ �׮�X�}E�#����d��g��,Dj�1M��I&T5�ƞ�x�[�l�{�p���)�9�)w��k(�:}��')��]EفJ]8�2�Q$��&��v������`���Mv�c�Q�[a�灛��-�q�u�@+�����auD�0YF��b1>Z*�� w���U�}���y�w�K���	��X� ����Q��-ŧh���7��
��{��II3��_�������y��'5�����]����ۛ�U�ʁ
8(�~�l2�㺅o`N��d��/WJ��o8K�V��D�&:�h�LxFq�H&�,1��7�ʱ��	c[Q�����N�iޓ�6�0�\��[�b��{�۔o��\��f܆%w*��]	����3^��l�ӧ��+�z��ᙷ)�
�f��Y�Y�yG�RO��D��W�`��ex�b|D'��򽬌��.�ߟ�]{O��@��#���\����Kt_���ˬ�J^@�K9k��� zĠr	���{����7Y�hJ6�^�>W�L1��֬�O@�W�l�OxP������I-B����-~��$η���P�V�����G����]J�����+��VX`)�"-w�і�eoh+����Hs|Ӊ+:v�bn#,t�ar<�E��w%�;��u����C˩M�MB8H9{�L�PQ�mQ<Tˊ`�<dG[c�t{)���t���Y|�1}�ﹿ�q� ����4u�$3�	��7_�Ye�"�Y��>���è|���c��e��e~���ɪ��B���_��Y�,��b8=.���10I�մa�����)���/���,Q�ཕ6��E����],�K���q#M�1��l$�ej�nN�o^�Ɖ����A,F�h��>�A�+���N�z|�]���V��T��t�����z��ܜ���}��������h^�������R|��S4�j�+�������#���)�\诖�,�Z6<www���6���	utw�`ea�x��3~�����U��T�O=L'�W��Z�()���K��ΣϪ}:�SlA"�6�I�B(�ڦ���k����IѺ��W��z�ۧ^�.�$4��[MbJԹ�הɦ������:�m�Ր�Ъo
1����$���Cki{�0ޠЍ�uژqd�Wc_q��l6��m��ʩ^�KX�c�'&�L�p���GN�h�S���g�'vǞ�x�1���D��]8Lb�֣6k��"�l��������NϜ��~`���ɿ(��%=�/�I_ѵa�#c�	�<*�}��8,���E�WK�?#�,,T�i��ж�J2��H�<��MF]���I��5c��ݢ�2���o��ud蹒x�$�օZ_�����MV1/�f#�(Ty�YA�\���)P�Z`a#�:�\��4�$|�c2��[����+�ed�S
�sZf�'�����}��a{�Q�dXsҴr�q���|q�r��ɝ�6��,�o�xgX�|I���W��p���2i|�q�~y:��p�v>�1�Ծ��V��zc�\D��==�(YY�_n�rZ�8�x�&f�%Ti��ڢ��m�B��}PO6�ݼÄ��X	�L��.�r��q���a�e�<�H�������E����'��kh�O%�|ű�%�9T���@*t���a9PL�9^)��uZ2
A��O2��G)�E� |��}f��h'  &��SGkT�G����]a���8��Wo2I�i��<T����q�!�:�����7ku �t��N��g
^%���v�J�_��k���`�O�]᭪Y�jqԼ���>5e	�O��v�p����Z�d�݌s��_Ί�(#5��J������j�7qN@|�īF��!i�ְ	n��y��)��}�����谟�Rs(����F�����:����9�h���N��x[��6�oHJ���ay�di��Q�}r���-�����t���,�Rn������|�a�_������oYq�vޏ���Xƹ"��n���<���q�HC���XzG;v�����p��ɍ��%�����h+���ez����^����@mڞ�T�F��8~Sd��{��y��'�:�:��}�t�io��+}#ֶa�/�@׼郿�^Kks~�q�8~1eM���Z�yE����;P
ן�8$+�8���ڍ?�k���<��"�~
M��w$U�G����P�&�d�˞;�%K�W�k��Z�]�3�<��*�\�K1,���	���@ )k��}����5�y\��Salf���(8�q�r4p��?�/���`űw][#��.{��~�*�ozs������b���T�"t�E�[�9��p!����D���d��ar�Rr��hA��1\�Z�����3�?-E?|�sxY	��%�"'h�ѡ"��p�bk����.���c�[Dh��C��63>�����Lԯ;D�#�cl>���|�*h`��bʉ�/�{�oz��d9��wc�� v��m�U�\ ~G'��V�M+� �#�@I�ۣ�#�����^q�kT�
�S��]��k_Sr�'i��p;��]���
�kjS��/�Gŷ\�<��k�<z�@<`l(�W��G�o�ʳ��䀊f�~U�X�|��Oo;�B0���_it%�o7b���Ꮵ�oj�Vޜs���*قa�f k�yP�aČ����� ��@���'��82��ށpc��g�/ѐ�g�s�x� _g��:*jHȼ>�#��Sč���&�a�/Z�mqe�A���L���x�5�ߟؾܤ��Z�����)��B �$X8te%��'W+&�R�X�e��I�ζS����I��H�+�e���K�D�lM�������rER�߹|?#�o�@ uFa5�c)��;O\�pB�sR�֔W!�.��+٪_(���*&���Z-H1�*���-���^ ����c�gt^|�����<��*ې��H.jt7\Hy��SVyU�������	�w$��X�����y� Al�ğ���D˨�:ː� r�Ӡ�9�9��nک�-��Y�Ř
48��&R��Qd䎖�9����^~��>!�SG�K�kWJ�?��J�/�K�-g��th_�o@�g�����d6����"�ml<�q%��W`�t�n�`�J��;-��G�q��+�C�$�1G����c�3У^©6���M֥1��N���9Ʋ�#d�\�d�մ�M:�M�Cs���vO�0��wue�7Y]r6o�I޿gBE�C�wZ×<���}q��P���@���Qi�ӎ��.4��e���y��L�pl2Ň$�(�p�*)�S��z,?m�쓃�v�:�wfg��A'gL����ׄ}��bmc�|m�e�#�5�g#i$!�ӻ�Ea�O� ���DI����
�d��s��y/��"o�{�'������=	���)��5�<���$G7]:�����=
ćA8��&!b��U�L�z�/(뷲�:8��F��NКjw~n��&9��d���k�r����S�g�O}�6����Η��QX���uO�^���Q�=�O����[n�s�\�;�'�j��1����/�&+(b�rO���#��^��Օ�[l��B���@�e��Q]���/=#��U8f���-3CÇ6V��c�d�#<���������X�;�;������|Z�Eٰ��ko�軜��=���������Ԣ�J�
z�����6�5�d� �93l� H_9� ��Y�����æ��+.!��+�ey��2s�2��0�]*�졅۹5g�OW��.9�!��}��g}7�ʑm.
��b�;d��n������%�D;�ӐLJY�p	�iم��e�L�A���ƥp�v#��ψ1N��@Zp�1B ��f�t:\!��ck4����5��(<|��;�gD�_�`��`^n
��i�5=�j��ۋ=n^�u���|�84Sb�����r����A=UGtĒF$�T�&���.�-��|HM��5�N%�fN���|���	�Ȳ�����OΌ�M"X�,66GtI
,X��[�NMGT���XPmq
�$y����_;!����1xV��9;��b�v�􏛸�4+�ٮ	qCHP2D^k�3�T2�ӛe�a9�[Ъj�GyT�[b�4�2a,���Lδ��V=���--.�|*d�?�i�s��������p]hc�y��n���.�[�{�	P���EDl�1���Qz�ǝ�S90�w�l��T[Ƙ4&��[���au��vj3]�S��I���(�}9�	�榆����I�9��v�c�L��=��T[F�b�B%S;?®�X��U��l�RG_�)��%@�#{i�3�&Nq�~?����{;�}i�7�_��n1���9�b
x�to��[�d�7��SQ�D��z��;�<�8��}�ށ	-D4Z[0���G,�B�7�ҦR�sl��p�0k팖�[uW��S"���ƘXz�vW�5ͭ�w׌��5�}>����e!JzQZ�~$�B��0�w1�ak_^��|3��v�6Aɗ^��n72x�o��:��ht�xg�>ȢO����?NkL�[9 '�.k=IHE�o�:��%�oC#�.��-�B~ۆ�QR����ƚ˽6C����qh����d�*��c���	���i1�y�@_Iڒ�[sz���V��|I�T_A�m+�yg�Q$S�׻��m�MT��L����xпL���ݝ��#���@�Qx!�s���<Z�vP
\�M��c��Yp��HzEn��\&�u+;��&����1�~t,9��X)�E�v����7Y̝ʔu�ܲ�F�9�Q�:EZ6i1�~��h��Gف"������8v��N��_8�"�c�v7�G\���!�N��u\�rs'p?&c.	�AMWnŞ���f�+K�1���A!�a�S����dpz��V#9(����K�D	����,-��^zeJ�Хm�K��v��6�e�s��t�x_�N�_T2������w�HQdd0;l89p)�U��*n8V#)"ڸx���^��C ��hq�5(V�]�K����GYMu���h�ѭ8tc�`zb�;5����5WK�����SQ-�i���q��w���P��Yh�B�G���T7���uǊ�H00#b
���s��zd����� t���L��蹇���;���Ij2HBkLiF"<�;�Db���zN�9�kl�������S�r����ꙣ&�~tL=C�4Z�~�M���r�����cEX�>����h%@�ۃ���鴍n�yo�>.�_1�ٿߩ��?�$����B�ӡ��&�q����
9K���qG�M�$a�w�2�7�������b��I�˃����WfD��2u2%�
��w-�RW}ň�xU����:��r�*%Ps���-��r���m�4/\���eKp�Q<��D��p���ƞ�9&�L�|�|��N��CHg ����BB��>�����M=+0������,���A��Ȯ��O+0��_�&�?�ݶqi��>�	��,NkK�Nm�����g'p�Fitɣ�S˶1��@3�p��`ǘ�U�d��T�Gؠ_�W���nb���#.*(-�k��3����j��#T�����1�ͬĂS]ʷ��h��Qy
VX������xą��*͗�}^A5�����`Q��ȤV�1���f�Mw%E�uQ�;�<�Fn����L�nV��J����I������+�J���	ʲ)w^.^���OL�������r�ȼb�N�������OPt`C?��9�Y؀���������WH��)��@o#'rЊ�������B���␿K\%W�ل�/��]B�k��I�|��#�Vp6�����ר�Mڟ�\���a8�Ii����
bq9�I�Tz�N��]�֒�O�����%�~��yZ6�n_���H��*��@�$�]�cM41pZ1�Q:WE�1Z���4\"D�<h.�dk�w�{\έ�\M>>2t��CQ�W +a�p�5�ߩ\c�6��4�P-�*��H����3���x	�/���C��aJ��b�D�A���@�))�lp�T�&��8Y�L#�˦��qRv�f1�] \K~�L����x�����TЃuRRz�*ޖ��EW��X�;���2���<���(�\F�,�y�*��� � }iuG�����`���:��<D*����g'|� s�`�6d��
� �+�1�;{]!I��jl�8j�:����
u���b�';�]*����Z�9�|&FE���@��A}S$U��\_�hB'#"$�©FZU�L��w���KҔ+����K��ȏ���t�Sy5Mz"���3)}p�����::T,����䉀���j�G`���W�¥�|�� ��%�+�P����T�MV��V2�t	�V ���ć���	��N����(�h�h���̢�T��ce�o�U�8�Ѐ[91�\�A�E�pA�5j(�:,s���0�����Q&<?���#MS|㩐F�����TE���?sӚ��rPHl���k�t���C��n>z���wo{�ΈJp��\I|d�щY�r�Z�U���������(����eR�^Nչ���x�r�)j� �8^��N���<�ο��2�K�0
>-v"(�E�k������@��^6ܙ˅[��n+��=A��-�w��8V�~G:��y�jKnH>���Ŷ�E{D؝Mj��N�[�>|L^9B��t�M,�n�	�E�g��=F"#����LĬ)pz�Z�2��,N9�y�#������$]Sm�YXK�ס��+.a�ZZ"�>m���-^���"�n�p����Lݯ�
��4�Hi�XHj�ggN�5���==#��%[+� v�/ ȗT�u I;� �٦O�5�7L��`0�>~v��~*��~Jj�Ka����@1B���i�i��:Y�ޖh���؅��x�Z*���9�I%�55R�j�up:�����y��k�� �A"Z"&�2�f�	������r5�컶���k��Ia�	Scl|�l=�An�.����:���	�0զ���D�ړZ�F1ŀ�ü�����b>�
���JEi��~%7����oq���P	���5�.{3��??	�\�Q����S��+6��D^���u���h�pw���X�� P��,�v�%����Ϥ���IS�r3Y�v��"Ɣ�����7�E�&�ԠRQ���8�i�v�@��-?�;��1x��W�8;@��t�y1%F�n�T{С*�ЌG�$���� q3�h�k���^8��	�`(�}W�O��K���?�*j�R̅ ��(�^��e�
������w*����#>�4��p.��a�ϋ�F�8O��(/��_4���] �Y�4����I�� X�
gd��V	�T#G���+B|s��1l�W� �t^�oZ-�XIr�l�Ty5A�җ���L��Sy����OM��4�'~��)�G�\3�_]��v�����\�q���h��&��me�������͵���J�!�#�,}�d̋n����ĒW1.*$� ��:"�޲���|��+��h���k�}�7o�x�ɴ�����ߦ����3��ۯ�^�è�cj��B�l��,A����[�ykK�#FF�m��u7B	��sډ�2rK��N��O�p&\��¼̽���M>�JJ���'��>��������s�4��7�P�4��D#3�{.TB@M��v��h��2v~���tD�"�k�2O�$Y������e�X��ylR3}2��L�?��y��X]�+E�?�a7x�JjC��Ġ���4��?_f�S�H�Su���� 5/h5��D���W+O1t11q�g�v1t���Igּ�D�j��U������։\� 3^DwK�*���45��=&��y�@�5Hp��)1�������_<��+7�x�K]%1�"M��W��yfE�<������_ N�~1���˓QRi���^W��`� �hƩ���:���A9ңn:��0��� ���A�}Ӂ �D�$�柌M"*lN��w��!�T�O��bD�Wb�!Ob,�8#o8w#����v�}+f<OB��� ���3�H���gܭv?��"pL�<�j������,���%�H�f�8������Њ��%�5�p^���J�Kc`ً�]➺eQF
�
����B�.q������#��#߿O��[ƥ�7����d N;���� ?�xVڑG��M�G`�����7�C�80��<T���.���ԝ���'�E�2R�)FX���v��]��_o`���ё,ů���	��-��;���X��b���"��wN��N�鼣W�a�`c땿8CdG�n����kē9�E,7in~�ʩ�������Z�����,k�G�ƵJ) T�3=�~�S3P��]����n������V���%�h��T9�V	Uc15��~��[���YfyM2�@�nr�YW�ƣ�ؑ���+@���H��vop��a�Z|���zɇ�bU�0�@���5�e�%.ya:IVڨb�5�6� 54^�KJ���pe;��&`��҂�@b6�.��� �@�~ю���=��ek�{l�kz�<��KSJ6<1��Ņ��C�y"
��9H�S�d!ys	�N?K1t	(M�곟e�փ�V	���F�{$�o	I�ޟ*%!��JC1:�9i6#F���|VZ����~�BH��3��k��{%��Xى�2`�,( �*%ր��Y'	��h����0��m,U_��쒌����E�u��0�����_e�m^Zڬ:=�L{���|��<�wL���I��F!�1��d>�($O-6m?�0+02��J��j��ܐ����*����F��}�]dJH��bǹi���Ŝ\�)�gY��#S�MMe;("��U�`V�29=���g�V��Xq) �c� Z�z�B���Wy��?��)�F�)~�T�0z�7`8��:;�����Ɏ�>|�g��!�}�?p5T�oj��:b �##��n:h�W�;�
�E*�����,ek�ֈ`�o^��Q�Qп1ڻ���JF���͜���hVG]���vG�{��D]# U�gΣ�0j.ә�ߥz��[���E�S��2�@�������5��!�=����L �2��Z϶D��� �$���!�� �a'�ݦH�]��*?����j	���>���@���*��ud��a��d�#~�UW�Y-5H��h�z{�����13!�W¼�|s�#4���E����.Iu�,gj���(v�4�_��lhUI#��[>��@�fʼ^��7�� �ß*v�m�~�8����q�a��Ф k���Q���(�ɪM�ֆO ����u������E)��n�H�eR��g��p�)a�� Gv����&9�)�����I)�fH���4�h���[�):��U����`;ŐO���Lp�*�Fą;��k�D>�RF�&S����ŝ�ş+����z�fpXC���Ll�$�ڷ�"G���966/�e8�&yHHO~�Gb��^���o��G;|�F6��t�P$C�<��Wyl�e�vR�^i.�g�c ��㭖���oﰵ��\X�U��J9�K�?���=vP̯����-)9��j��ئ��e4v:�g]�O�Mqd1�W�w�ur_��v<�B𝵜���;�Xrg��\���j��ω��;���=����V%�ej�:��������f`c��,M�y�YG2>W��}�PT�M-�lgy��s��\;l�Ou��X�*"�O���;g��''�� }$\[K�!g�Y_| ԾG7�g��A����+�,m/�큙��4l���)dU���%�Xw�"��:��W%)��-O���s���R+� o�u-8vY�
)��)erGF�����d� e޻�rƌ��h�M�R��`�Ϭ��~�е�PucːX3� ��a������e��xr&+��נ8Ͽ`�ʪi��f�φ�]��I/�Y���u�%��|:��T��p��,^B'���s��y��6�r��24�,}t����B�ο����î��2�# �e;9���(�Y�������qi���ݞ�|�K��v��BԚ�P���a�?�B @�4C�%D�N�4*���� y6=��@A��h�(��5w���B�7LF������Qӽ��>~N54����i]��t|M����m�W��XP&n�!����EV�ʍ�F�SE]\��?��«<�ɺL���X�M��K։�d��p�����t�;���w, T��"ux�p�z�~�^�R�o9��e�&(U��5�|'��#Z߽�*��7C�"�u5Sޠ�Eٞ���ciobUh3K��-�ch=�BwU`̖O*�6�}�s�=Q1�W4�a�^�X�g�����s��sϦc�4����3i�� O(0x��aص����5tWu�'����UT��;����Y���'���5��W�ON��;�Ql��)�$�gc�;͸Y�L"�-�T[�!�o�����<躼��k�G�����3�PN)r�zfm�3J���FG��Vt����7o�Cb(����mf٧�Z��qe�bh/��8�@|S7!�Tr8YE��%��������5N����Ϙdd���	MX�������(g��V�`��Rt�gw�y��:��{`3BA��U�e޹�i�����~�ϵn��nN.ֱ����=�������V`�8&�X���S�eqr<���T@j������Խ,�0,�]ϮǴO���	�4�T��!7N@1��T�yݥU�|�����\��$�A1��«��.v��"����{�$e΃�F2.N����W�Ы��5���5��2��ط��ZV�j�Ȇ��W�~�TIXC�V�'g � ^Dq8g
8�\c�d̜�_J��w-S$_g��qm��u���O��&�9�pE3��S�D�94M�Y����-n�"�Bۥ���"10��2��~�N���J�  ~��� ������%�v���$-7}��JV�����P�jt�����U�
��ξ㝇�4L����}!�4�Xzb�66Mv��+���ʬ��Jd.�Zx52��Аm�Ĥ)�&�;f-�+m�+~�>����;��CevC�A����+}f��lx���IR�9j�q,s�ڡ���BС�ǋJ�����~n�蓶e^]������a�Jx��hP�_����c���![$����ڒ�ۦ2�^n��f���цn�����9����%��m��t��k���f��E2����j�M�Gc6�=�MM
�W�7L�g�s�e���:B7c,<�'Ϗ�Ue�}�^��&,�v('�]�\��s,�~��sB�[�Q�px���/ Z�$|�n<A!O1;��}� ���3���Vq̫yj�՛Y"��/~�^��b����_�c(���
�v���3��|U0�����@>N��1m���#��Xc���]O2ҝ�RA�g",��PَBV��G���/';jE����'�g�`bȪ�[�e�Ӂ,�,��Q�GV{6�.�k�f�13 ;��!7�F�y:z��'�D�ӌ��sz�Cc1z�2{S�ݟ�!�
n��cܬ$f-Ox�aԣ+8|�i�7��z���'���7�3����m�'(��u�. �h1	�ԧ���E��ۥ»�!�Y�(��IV��Y�\��CkTQAʦoc���W�1�f��[��$X1U^-~j8y�|CYG�7	8�r�Yέ�(�~n�C�UG���I�%�C���!@�஋��[ �;�Y�=,�����6�ݽ����73��տ���n�mA��G�`��F�sC�+�V�1Fa�kX�=,p�XL��;h�1�#[�����Liy���kܳ�TțSR���v�~�Hy��l��E'ʭJ�4᝵�=�ș�ƒ<D}��B��~	NY�b �n�{��ɹAg	O���p�a7S;�ώ�rL�{�:U���
���Iw6i��5�t� �W��ʓ�̣1en�~� ��z��NUj��h&�\׺}�^�h�O��$|V�9�Q'nAj�җ�%;���^��n��<d�~F^��_�m�"��@yq�ԫ1SuK�x��,�4(�w��=�?}>�Av�tln :SÓ��9z66����] �֮A�������7���#�U�'���H
�{II�ݵ�DCG���	t�������-X]^W�r�H�є��1�1B�: �5,����q��wO�����S��%T!�J�sj�=�"��Q1/1��"��V褢#�@������H��TT1?���-�#��MC�1J18β[3���'�ʄX����Ӵ?<�^M���-�_�����ȷE��H�f�-���cL��;�]^�ޫO�;`h���Y����RҴ[v�;{��k�/�v��;��,-݂�,)0�~_���3���y������a�-<�v��t��S��?�[B���2ǟ���ba0Q"���I	>�^g��Y��T�^L�������{�� �[4��	�1q6X�!�K��d`|��iZcc�+���xm
@M	LϪ��|'�z��K��_�q��eE�~k�Y���û^��S�,�=���e�rji$�=�ZL� �s=U��
j����������	-�z�^# :d�g� #k���5���1f��'1Se�R��K΍����_ۢ:j�k��b��u���T�zW;����O�����I¿�����ThE�� 8%{ٯ�Ro�n:��4�w�)'��шZ�(���G���TeǢǌ�8H:�����	X"�*f��O�V1lg]��8=H�� ��y'�yF�7�V�X]Y/N�$V�3�e������
�+B�l��p���X�R��#?#c#28��N>��B��Er�>#�U��җM����O}l"^�HqJ�e"!RDX($��;U�bO�'�������=�x���.�K\��Gm�0�@���f,.ƽ8�c�X�UŚ���9�zp�Q��IF|�Dm����M�̦����'�݉�/�ˎ�-��-�P2����0�M�>�A*���Φp�~�`W��s�0��aΩ�O���7:��u2��(��Uy1�ǎ�Q�d��\~?o��5XwM��G}�lHIK��� �1������Aϔ<�������WsU���{\QP�)
�K�eґ��O���?�$��i�-
^��ܘ4&���c͆�U�E�=s�I��D�4� �B�����r����k�YԢ�H��BcE��,�QԾ�믳1���.߭ �󍖐4��'���d�/5��=$6H"ܜ��,xP
z	�k�=��{��_]*�� ��J�/�i�H����6��V��v���qGP0��&�������T�8�c���w�pCq �%OhH\��2U�&�&�s�:Ҡ����ʲ?�)�;����$!|3OzE�h�p7Qd��x��&�p.���� ����+�82�}��-��D�j��/O��QQ�VXzb���@�N`��v��K�wˤ�1f�5��ԤR$N�����"���]Ku�+�d� {>ſ�C�ã��T>�@�0A�2��r�'�Mx�_��c�RZ-AFh��yJ�G�p� %<�X�R˫ǿmqڍ��u�8POO�9ɗk�b�	�<��BX��z��7�L� �O=����zY1�}>$z<�̈́�״$$��^�M< ����K�6A%,<�:Q\|F�ǯhM,ۏ���^# 5��:ƒ�iǔ+�Źh3���Bk,���/��aj /��M��j8�4R�[�I�7�v�Ǒ&��cC�{}uBiT�Ɣf���]"OA�Q����s:���Ǫg��A�<�i�qcMt.�#s�G�e4w��uhEIg�� pa�p��q
�<�)X��p�Ut(�}34�q\U7wf�/**��G�5�P��$ȭ�0`8֧P;���4$M���4Kי�bZ�"��-�9����<�?�~�\�*��N��7o���>/��l�-�J����Q(;4^[�vQ�<�Ne�_������S��(*Zj̰d:@L��!��������b\o�_Y�(����X_̡,*
(��Q��ZQ���Ґ�V��ef�C��6�a*�Du�����MJɶNG��QNƞ�:�L�#.H���M�V
���H<�T�2�)��ss���<��<A3���k�Eϭ[6M�v�[�z�ׄ.��
E5{Ppy�Ǫ2d�7E?&�f�^�9�֥4�Jp�� �HMkA<q�Ê]x�6LZXHL�4R[i�j��_���Kw��3�(OK�t���k�^g�	Q�� ��O�1F؛�P$�T ��IE��O�f���$�Z�%;�u Oi�t��b�3Pg��{��!�@��غ47���g��c*P�(�+��UtEǰɶG��[�b�t���D��3�<���3
.�j��%\���� �ݙ�� 霘�ȑ�vcM�[/�+�I�*;�:��\إi��$��wAF)>�:��9$��$�'��<�U!,����p����b��}gw,�{��= ����$��w*�|��?����U�>Uq����G�[�L������(�P�xi,�Hd��
��3�X�q���������8&�0�F-0U�z^/u���i3Ai�I���%
0_ 9��(`�DHfɤ+,�ڣyT������<,�k��K�(+ ��j����OBfT�$?�|����4��7��^T�@B�Pgr ��!V�\K���ff�)=��EԊC��1>?t�>��m�2(':��.n��͒�Φ^n�ޠ�~��d���� :X��Ȥ�FK݅�Q{q��Ɵ�HE�����u�g�k��X�^l�%]��n2H�Ӑ�	�h�
}!v~�"=5<�+w�+*v�JU�V-�e&��/�M��mM�~���K������������WǶ����d����V̍����\��]���'0��l�!5�a�=V�}���=hʢ^�#��lMIelX!����y,Ws	>��Zt�8~���~�F��7�za[y�Vر9Y���شqf�3��>*��;��(v�W]��L#�W$����A�|�!�z�q��{�n�w�iQ&\{X�+"\�	ڿ"� {�����ѳ0W���W�Q7�h���"�k������˯H�IWWx������9!�w�H3���C3 ��1�d�7��n��e�ˮKk~ؕ� �i�.�3'ռ��#�)C����|��]����̥���|;��	A��j'�I9՞�dpty�n���>�#���ư��K%��T�
�˗2l�ߥ�}��W}���
oP� �������抋����ÿ�_�01a���=��6�JM�u��>�ul6��N/(���sPF��	.�M�fdi��]"�����kĽC}S���d�-M[�$]g_�n��+�1��b��'Bm�ú�s�t��o��}�	�[��|��k��OC�"$�����d�%`���k�ޮ�-ʞw$꘨D��8�?���Λ���,~F�EY�z��7���va3/�k�h=�il��U���y�ʀ�
�@IՉMVxCyH���8v�r2j=�Й8k�u)�-͋�$O��j�J*��4��S[�fc�r4��f����򣀅ILľk@�9O#�B��s����RNDk�Ou���G~�6���V���i��u�d���#ɼ ���i�������w�|>�ŜÝ�KL;?J�7eX���H���N7��S)є�J,�(���:�>EO_W\/�[�!��~�s{����]�$7�%������OA�́�~����p{&�''���[�;L+R\.x�d�{]u��n��WXa+�G�0��rO��ȴa����B��7��G
g\D�Ie`�+Xr�^�5�L�$h�i4�RG�Jb�'�m��Ґ���5�ێa|�!�(h�3��W�2�Zu��;�NAPN7e!�b(�!~'ϱC��^��ݼ��e-����+xrT8��޹q�t0�5�F��믴�6�,P~��U>yve2�NJ��LN��3�S�A!�}�"Z��|��ů���/"P��0�$�0�Xiowc^���<��z�q__�c )	/��$#�3�[[%aP�Z���T����\��7J��N��8�9��\������5�fo��SWB��2�,ԚE
���0B�֍�j��v��]�]�2�/�k
#F�X�?%"վx�G�^��_ȓ�R[����`BF�����������r� �����:QZt�PW7��B�o��.6�V�Ii��!]r"��r�=<
k�1xQ@�����Wҥ���ש�6��p��GL21o�%W��y=$��^�T�P�w6��B�H�+~Y���<��G'����=��'��q6W)U_h���c�P���YrK����>�7�U�'Z��I>�oi@r[z;�so��)S���P��z��A��<6���%���5	�뺰�#�����4u�/�77�|�������r��8`�1�7C�Z�d\�~0H�b~��:�����tGվ>hE ��j��y�N�`ⱗ��Ղ�BӞ�c<Ɨ�P';;�߳l�w�gڒ�::��=����l+T��%���I��o��ӱ�3S>

.P�@��-��`i��n%TV}���a�<���x3 ���ev~I7�`aPכ�Iw��j踹T���	�%�k��|u�,i#�O��vZս�nE�Gc�<O�w�%6�3}� G�BXXkQ��;�ĕ�O�'�X0�cx��f�G��Ƨ�$S�jL���O�\Q��QNP�efD���ٶ�"fpUR�+����k���S�n�/O�Ԛ�`d��`����X.];�ɮM�!�E��$��&�4=�	���g��;�(9��;�C�6�؛��!��οMn�^d�����y�Ɲ��pP	2V'~L�8�\<U��M�G���Z�uI� ����Q0EIXV̀�o'�\��o����=�������:;���Z
nٺ��XQ_ڰiU�w�t��ӔH�w�,��ਢf]����>���h������:�0����U�Z[-b����Ji���ءQ(:�����:v:�A "	������䐿��5HP��G��CcK,b���Pݭ��|�v_�ua;3�/>?+Z������N߇T�y�K6��x�l�����C9���t�[�ɉ��t��TFWhմL7o�Gh��h-7aPل$!���g1�`�f
 ��l�g��Q��P/i`��q!&k�vmc���<�s&�}��ޝjp�?@`��|A�n��D�J���$��w�g�.�2w=�5����B��v�����R7n�RrT|�u1�>��nQ�B$L&��)M�����l�Tt9�������P�t���;��dh�\������>�&ĥo���:��&F��cB��Z���'��`�}}����i��D���6��U��ֺ0"�&����]���V�M���-~�����u�7i �U߉���@�bG��	�8�K&�� �>V��fiHr�P�ݭ���&��[hj�a���x)���;�e� �����y�=e�P��Y���<o�**��n��l5�����'xU���䧧�Z�ea��8l!��	��Yrg�~�_w�<:��ʑ����'�|�כ�F�<FM�i��7+��fG�|I���F�tQ������D��n��)`���ם��ӪJ�����zbP��Nᨶ��%}D(��I���GU돢`��n���� Зc~��_�NH�D�$%A����
�k�[+镟����.l��j0��ӷZ �n��H��5>�9wx�+E��'���I�G�+2��&~X�}���k�s�d����$I�<��ڹ�t�����!>Mh{SS���<��!���-��0�����5��H�1{�/����0NKhY�$94kӘ/[]Y/$�\N֘�,@�}N��ኁ�pqׅK��K����������M�#3�vf�������:���N�����YQ���k�)�su�K�"%xAE�Z^I�!q,�S4��,.e���ްc*ZnV�Y*�{���� Je���<�7�y�����bZzWW<b���Z��%�0��k�Z�}I�Ϛ��ݽ��b^p����\��9���va���~�_��E|���!���T�jN5Χdi"$�(QtЦ[#�ը�$��*���nB��b��Q�� ј��"�OY�Kڠi)�f)�<�5=��C�B�6���}c��9E�a����������-�P¬gH�A�#��F��*�;c/�P�ƈ�/ d�n9��x4T�	
$ҔU��BS��0�W�YB�mZV����*A޺���ŅO����	B �zY �Q�*	�����nD�1��4����bɹ�a��,͆S�9)A��@���:$����!���o`6ږ"Q��+`�
��A�Ͷ��4s�����9�=b�$�L��B�^��?�d/��Y��o�f)@$oOK��%����<U͉y�����������="D��jַ�L����~l�Մάcg�����7J��"���V��B՜�h�G4t@1YVݨ�N��E��h��HM���kε<��{���)��N����u2;WX�k�b�UQk�-�L�����UU�73��z���N ����A�S2b���d{՚��Z��w�w��JN�s��\�kEZ����c�ZzI(��8�|�ilY��b,U(�U�B��5аB���f��gi�:Eaϧ&s�6_�k�.���k�����ĳIF1e��Bce�lxa�u�����>B�}8y݀v��bD�
!�����@���xς�q��R OT��/p?nc���@�q�3ꀢ����((:����J^&���]��ڃW��Gy�;G�4�h�eG�.j�3x�@I��(���GR���w�/������{��j_�f��� �������
�?4˔��bz#bz��^1*y(50��t�E��e�/iY4���!���0C^��v4��[�!%mdD9��>�b+���`��-��(2�zv�}�d��tk`U�'2-��ɨ����������H���s������D��e%�����N�$�z9��a!�Cv4}|o&��(9����^�_���pJ�����>C�Y�G���HB�* �(��L=b�G4���El�za��]x���5B����.�G(�Q"���&����%�
�o+㪫'.�R$��!��1�\��<ᯢY���ɓ��"�쬢����bjjC�Z�ܗ��%�}̬��a���V����u0%����i��?�@ ��6�UV���UZ¸���M�*�u��3:G�@�ڝɑ�l����I�	�� �ø=뇢fA���>x�N &�.�����Wʪ3�FJ*%Ĭ�`r����!=�`�O@�}���5=�r��%���-mxqn��ɶfw�jU)EUU�߽
� ��K+	>3�����^jp��\�)!�4PK���lmݶO�b�'/(2�oA7 ��(h���@A;#�Y��QH��h�_��*���A�������A֫��,���b�g�_���gH�i�GIh�xgx��v�kue�=$J��U�����#�HP(r�7�\@3H~���8k�I.8��C_
��ȬW⩍E�l]XL���r�^Q�XT�#6�C�gq��s��Ф���w��,�0a��_�F��	6m[0��$��p��-���W��GZ�rn�N/�6㋏���_�����ky��������xPLLp}�QN	*W�'JG.Y����I�Qn��rk��[�N�0C���OVk}=��?CUF�,��bI��#6Y�����ʑ�RI�Rzk7Yi����V��a'�2�K�����I��Q�|p��*4wK�C[[7h�NʝV�U�8��:u<7ΗD���=��}�W׈V��ʏ*�����1-�u�lc��s`�o���ܿ��Z6 _�=���
��LE�$�m�D��R��^���s�,�
y����M�-��.f�Y�B�
����&A����P���T�u�ȁ֢���'<ߛ*W�!'[���)��O���BBsz�m�#�5<���RS�qQ� �@�4	K���E@W�wҟ��F������甆��q�J��pp�?�4�����х�Z�a���|����Z5�[�`_�,4��Rʊ!!h�$��Я1���I\��1���l+�ܡ���p��g�&�o.re��l22H�[:P�s>/^�Ό�����V����ݮ
�<C�z�' Ϙn'��*��8�/-�Yk�\�}DqqP�AO	�Yn�nTA�*��K�^N��qe�U��E��7���m��%���s5x����g�}R6�������IA�2V7��_�FFPX���Wu�_�xㅱT6�ڈI{:�SrG��/�]�lW�km�V�:�A��P1�>w��ZB��	)7�:Gz�CpK�+B+X�$�7��&R���<�֋m��&r
^8t�I~��[¹���f����-*�Y��_ ���0RK��#�J_�+x���h�a~��u��3�`̏	/B� �a�v���3�pp�UqؕO��e��A�\p;)B��ٮi'%�8_�rI>!M6B��䖓U9\W2�G"8��w�:7������9��zbj߳ɣ�sY��0N�ǩY�:�
�O5����t��X�=(�o�:�5�N��x3��*e���$5V��Y�T9��"�����#��i|z8^o'k��xz�����n���rډ���q�zPD�oP�l����L������İknN���K��5�ꦡ[؀`�#:b��.&��h�>�J���k~�՝E}�T%�C�?s���'�!����H�搑'kj�7��������P��}�C�3��f�tyH5�Hqd����l\/�Y����=!�1�%�$���w�̀���]�B���u�������Ol�t;�9"�^����?��P�^kXİ�I�8���'t���-�-��U޸}d ��d�usA�Rv�Z�3�t�Eã���.���v'��Qpe�99
彊o@ �hr]�MI�&OV"dC)��ŃbB��s�v�m�ⴝ{*�K��zb�^)�V�����2�A/��(>>��������#�����k0L�!�Ф�B7'S�H�W2��;��,C�}�#�@O��A�(�j_eP1!�4�s�h1�� }�����]�X)�3d@L�p~g��lx-P8d��y��z�:m���T��Pշ����i��l�R�=X�*64<f1��y酩˪��5P��k^�@��8xII?�~�T+�t�>�A'�Ҩ��f�F�He��d���ү
L��Ʃ�5[.��Ku���U_�iO�~T��mרz�	�,������
��ܹӬo@�iJ��o&	�pfw�@��U���l�T"��c���be]�k��KCWN󉱨H�ެ&�۰�L'):z0&/�+����r#q�(�A֯Y�T߳&F1q����Z�T�9��e��;���DY��J�[���O"�;Y�K���f49�q�&$��t)ATl8QSRc�Ǵ��X���b�#L�a'�&a㵖2܌�%��	��12I�q��m��c�_%3�;7�P��U��uw~�a������Ƨe�����;�O�����2�H����4��VW*9u}s#TW�N��伍��F%������TQQe�V��_5��/���M\��{G�K?�OZ^��qW=��A�F���V�����<UV���M��V��7MVZ]���bn`�F$J^�����-УV���K�w$B)f��ǁv�d�9JU��Ro�g��劸H�]\�����5rTP��x�������IB*zV�~�}ߪ��ȀF^D�o���J^y�x��	�Cb�۹C$���'L��Pnj�Y�k-���ܭ���0��sG
nj۹:�Y��HB�;�N�f����_�������j#��}��g~<Ӥ���꼃�C*vv���)�P��*��kw/Ff�l�f�9{��yoդo���9��ȓ<���d�9PH�������[:gp[׏�:}�Q�t��Q�
���V�)gP����^l���ɺ�r���8�!��?6�+�f�R���M FIϊ���S=�����]o�׮��NFQUFN]�O��3��O҂� ��9{���ܗ��#��N��_����ԕ5�UU>Y�R��OV�U"&U%d�'%����լ:Z�{ܛQZE7Ng�?�^q�Dko���#���OU�����cG�a�w���I�>�J	���Q��Č�����k1��F��V֋�L���_������o%��jL|��'����w�j�u��%"�=�̏=��Z!i���LQ�IYsk��;p!:������%u������ڸ�deӴg���Q>⊾�?hֹ�ۢ�[(ΏքU	����^4
�%�E���X�/j8^��"y��<�>@a�h�޻����9<K=+&���H����i��^�3U��%�|K0*�t��՝.��|'9�Wi	y.c�W����F�\�H{�*ص���aϳ��6E�*��ST72�,8
+[al2��j��Z��6\D��l��<������}ԥ��(�q���B�ίG�ǅm����[������7�c+4�*Z�m�Y�Y��=A����u���q�b��� O����\y��<��\0���^s����U6�<%�
ծn�ѷ�m�y��H͈h�ަ��b+쪕������A96�ps�/*�5(�o{���f�4)ag����o�2�`��n��*��`K_�ő�}�(6�2�Y��m�̓�����.�Oa.0��/5,D/��#\�Z�^�VUx�fw�{����xt�W���?�hV�<VoY�Ԋ��u��^���;UJ��%\1�����\-?OM}��W���*�9�:�SPL4_��ef���a�E���G0x�S�ʲ��+j�ۗ����wQ���ڇ���Ƀ���zh,uY�&��C��?�p�x�0��~Mu�����N�Ш^x�
���׮>~g��U�����N�u+/����B=\Z�( ���m^j���7AZt+l��D<0�X��B+�Z�\�*�������U�V?V�)�.6,��$^?E�iF�5�k��.�)*~8®ҷ���C/kfl�E�e'�,Ƹ;*r���u�lى�߄Jޤ�t���r�?�0M�W�������� {�qV�'�$���$R�<�c�;
�#=/�ݎ����� ͵<Ά~���Mz�P�2S����1X��Ē��)��W�iW�TŔ�_����@�2h3��� ��Ơ�e3�P
�W�	df#d'!!�֟�2Zb����m�_6y5��/\R
�鐞'�掩�<������Y$���v��Z�ɣMl�M�Uv<O��/�l���{����ĐO�*�	�F�Ȟ8ב��׻�)J�6@�S8�V���6#U/��ߙ/�}l�("�'��Td�uw��>���ֈ�8���6�4�ij���A�=^��7����?_��,:�G���~�p�4�햊�MO3l_��_�=?5L�M��i���:=D���i�����Ce��mˣ�]@������6Cص��jQrb�t���� zl��ܮ��`�����N���]"%��m��o���7+|ww�A�Oڍ����������l	����ދ��t�́X2ݟ���v�����1�HVF5��}�h�IV�
Z+�ْ�)2�y��3Et�}5&���ug6hI^��le�w^���Ż���ɬ�C�4q����LH��	x�j^Ș l)㆖в-=�>>����ј�X�v���0~t����]�S;�}H��Lu�"e�25��������z�a�K/�a{���2~�b⭳'ݵk'�Y/�Ζ#��iW�~���XY�Ol�_n������VEr�u�4�φ�})��Y���#����?���'2?2��ה�..&�g�.�}�'M!��JJ�挈�n���Z����
ɜ��<��EIc���6xH�T����O5G��.&�qde�wU�����t&��*5ORy�vǸ��|�hG��#��&ufp	����P0��v3�����@�ҭK7lg'�S�x��]8zj(��լ�.�Ji�:\�3|�c8k����:w�YP �F?�������0�̳ޗǛz������Ԑ��{�K�1|T���g�N�uV�4�:��o֗#O���,�)�)Tl,�ɺ^78�#�л�
ac*h����ԗ���������W���	%��-��ާHt�K���8MkFz9�O��tc5��E�|�~��$�n}%�_݅���r�Y?L�h�3Cp%��X/����*.hg�����6�sJ�	ˠ)��E�S(55R}3}�)ܗ��ݒ�޼�g�Wpۿ���
�i�>S���d��0<�D��D;_I���!Wm����b�=b6[�|�?��E�w�ob��[]���k^(ao[N}��އ�쇂��]�Q�������ح�ZT�������nQ���Y���]8�*���|F%!r�]ZA(����..יx���s��?LN�Y:/�q�<����0�G���pI��
G�K�=I��z(&0�<�r��|�K�5�#��݋A2�ۖϦ�{�FN���nUe+PkY"��1n�E��Yv��A�m��v�S����tJ]��g���x���O8gu�����g��z�i,��n@�H�uu���d"^?˓��L�>H{đ2�Fљ0H�b�?�+鲧e�^����6�>�ʁ���5�C��Q�O������%�(C�Qwn;v�s{w;�������;�L���4/��<> >��շ�vV|W�/�����uVI>=�.��ݠi������&�����_�}ܳ���xּv=���y�P�3�)�_�utl���9����}r�����
\q?7�?
�d�=��"MX�2����7��k#�����W������G}��	i/T�*t���F��`%��1Ϳ�D�Ae2��o/�aL����]��4BH���M�;�*ڠ7:��h}����7��ǜ1⥮��$V}>_�Z�rV{�����;Q���U�ϛ�ovkoL;p�cc��u�����ɴ�tnq��g�@�f��iN��{���&䁡H���\\|�	N������w;�L(����zԶ�3�߅|�=Z��6���[���L��v�U�k:�9��ddvf�K	��/	R�"�y5��gN��*
���|��t�L��|t�y}'j��5�jv��M
�[#b ��>�<g8��h8w���]ڪδ�_>�HJ�P�ɒ'�q����j86��2��B�����zw����A�i�䰬!Ę�C�gK�k^�醴��~�Je�O���^��$�����M�G�X@�{��i�}Ӊ�q���77�w�wsr�����'�:u������Ȧ�j�j�ֿ�~y��ׄ�5Ѩ��@�a�#`ޥ�?�[zF8��A¤[>���V^��d��2�\O���}���|Q���#�3�u?H�ml8�c��H7R��E]�$�ْ�͖�c1X��oƚsm�2��J;���_�H�U������u���4Gm�3{_�m]p�¸��h�]키=���9��f�7��!!��.��N7�ޢs��H�5��� �Z3�6c�f)T������w,�ұ���Q�p�f��Ç��k ��pw��#�=̲�'�C�&%I��
W�] �m0����������0������׮Uv5��PZ,�9�;f_�V��Ҋ��"��ٱ�*�i��t*U�C��&�Z9\���:�1)%"���2fM���K����ӝ��0���(�z����Kh(��y[X�zJ���8i#8~�J	��dG�&�[jaV�����sN��u+�0L\xx
G��#�R��ۅ_���������pE�g����Ƴ�j|C��?��L'IIǌw��Q����T�v����fL�<"٪ρ���1�R)�Uf�k�i_���s-����녖KN�~��@�3v�����4y�w�ηa��w�x��^kX'=�(<>�k��
ЕFi�|�[������b�܆��~'�NQp�m\�ۛ��������	���#�E!��Hg����qа3�G�� ��3��	��)K.����dO��?����>�]E�^m}F���,z
�h0Û���i��r��RE���a���ڿO��:�1�Y��C���kLbb��O�AQ��"��q-���﯇�B�������5*�|�,rh��2�$מ7�,
�TL�.�#�T?ݧ2�K"WT�ɥ���E��~���9IvQ�sm0���"`�Jd�D��a؛j�M�%��
>�;�<�����W����t�������<��L��D�N����$r피�����"��|π��U����>�#1�D�~i��� ��64j��@y��<P�6$y�gDFD�cd�}�A�D�q 34�b�͆ �����5�,��kl�΅6oy��{x��ޟ�,3�~@Ŕ�WTi�&�.[�I�I������p���-ݜ���Yo��_3d���m�����a���=���Ԯ-��khd@\�`�9�?X�9�ݏs83�-��*g�|���5����NO���>��ǓA�Zfݭ����J�T5IZ������h����.`�����Q���ӯCy�3�aHv��TJ{���Ŋ�g���$�	C$�eΧb�`�,kF0x�Φ����/cȋ��^���v�dM��\(��{�JE=�'��ML�w���q𙧋��v��<�rU�`�0]��&5�k&�-hh�#a�1�R�=���ľN��#��1�4IRp=>�Щ��da�AGA���FAh��v%?R�=��(W���/��t]�6�QA�W�$%x���x�v�w-��U��y�α9mh"��tHܛao�y���rBFF�g47�a��Ί���FtDE�2rP*��OZB�b�hQ�S�q$����ř\�m/��L��ڣ(eҸiʜ����.�<c#(X����/���dM�?(�ۭ���m��,�y�D�C���)%�#G]�А�����f,��y�;21�)��o�յ����M�X�|*+ �V�ޘ��e�T"��6��>ж�D������mf?3������g6�8�>���`X��|N0�%��p���A�M���v0;�]&�����5ʴ��*�vh�~U�Xs� )�E�;y���2�y��<��03?��-U�l �V%I��M�т� l�����(�1ޭ>�q2�iup�!�چ��տo����
���������s�� ��/5q�O'��4J������{,+Mc�����.�� b��e�ӭ���v��U�~"|޽fN�S�=7LD�p�x��bU�牖wխù��ܹc�Nާ���V �FO�C�y�_�߹,̝��~ް��|��x72u��gS1:I�2���U�ɾ��V�'�a\�E8)Y�pa�� ��/[EH�{ŝoW�#��A@��!���}��\�?�,bsv�'E��;5Y'���AjMB��ٱ��}���ڀ��(�&I=g�Y���00�
EL-٨j���� k�gu��W'�ZF���es$����1���񶈙(�J�9s�|F�9����T�8］1ö��3H�<[(�/\�u�+3O��7�����N["4[?d�iG�tY��9�u�eHR}�<��ANj���kx�0��߮�A��Z,
r��]U�?�Ҍn�ྵU�y3�'��!�
7����<���k	��yӶr�^���,pf[5�ɾMwCM;ؗ�'����r�DG�4�,��FTa[j�w��C[$�~�}����Bh�Z��xZ�B�{7�����!A��ے
0�8a��	�wk�ZwY�pt����\�'�q���jc����^�l��q�=LI�r6&�l��U��m���}s/2D������#�x����_�J��)��eB���Pd$z������LA�``�<��dm�.W�eg��Lo�BË�!b֩�e��e������`�t��dV�a#O���7�����^1ۭD�wf�⩬�M�l���9�s�ejJ��/~���-����v!ܶ���g G�.Wh�T����1��Nd5�4 ��C&8�$����<�?��~��c����튠��q��z�A�?7o�~X������y�S��5^��5j94?���!A��H�x�y��9w��4ߏ|�8�m�Y��k�`���C�{�@�9Z�V���ND)��Utث�4�"���A���KurcW��"�ǎ���!�����A��wϨ&��mto�(
J�ҕ* �H��k Q)�$�((E�7�i��$"�{�B3���y���9������^k�9�ٮ����ccS,�=2� ��Q��%��6��4z�	�Y�/�@a�:��&Fe�����˦���IV�I�m�	X����:c�*N=��}�\fR�SU��s���������N�B�HӀ�������^�ݥ`YO)W�J��Jƕ��P�ck�i�싼���k�˷ێ��B�S��8(��+Y+[\t"**����i)xkjKߔc��NIIXb�y�����_�y�w��3.t���ߋ$�z��$3��]��߀^M�!p�ѨP�lw�I$�b�\�hea���2��y"0UUqO�2�������ģN��m��l�z�\��#~������ȭ�9�"��C��!��~���b��7�#���������?R�彜�n��BI��<[m��D�t�ew�橬55�++�����[�u�r�ydG_�%�Flp�F�oae�a��cv ��Y���A��	^�6p�*U��(��hr�� ED�;0��v�"t�bu�٤.�P�<K�p��Ի�yjV�?oy�AZ�
��7��Q�x��|���a������R��ya:!��/��P0֒�k���8�Z��}�!ٻ�
��ίn��PT��!�!�Β��d��#-��op���y�,�yb"�}�Z��Y�K��8z�tW�ɖ��_�bS���@v>�-���~�;A����q�w2	'zRK�����侟 �j����V�q8�]�-���<fK9N��ۯi|���X^(ht>ġ�	�YMs>�����qW�,r���X�t�������@f&cS4�	5�w����yz�Lq�9%�-����D۬�`�jբ/x�_n�&?���MaD'��=��0�88E�d��F�=j�l���u��V�Hw���¯{B�pd��	��C��֜Q���<����6u�^C���ϥ�_d�S^�[���_H9߬��/y�j��YX侩�5�����Rb�|�FoݙF{ =�]�������WS���j6G-Y�%���-0�߀٣ʸ��NE��^^�:{�g){����'�1[���xr�,_g�`�@���qII����O�h�CŭM�)�F|���+���XWdՆPw��ǎ��8�Y1�d,}��ֽ��Ȭ"���'�2[ʧ��ʟ������ݵ���Cנr,g�_�- ����93ߓ�I�t����=��t��������_~'��/h}jc����%t�c--ޗ߹�U�i�(aJ��@�3��>T:P|*���)6�#4�?̏Y{��qE�f�-�ԉt����ͱ���jгr��?]&�@�|�u`����-.��)��M���� D�o�#+T|��N�J�T�i�'��3����?�I�Jw���TDn����g���
XU���:8
F��/��B�߅N�B��R��j���$^���4rB2g.�w(8V� 2��{�q���X��s>/��6+ujm��AW����f�A�Q�����G˩��Gy[�5�-�f^��ӵ"2[^BA��OvFi�S�E�����x�Ȁpaoy0t����y`f\3m�{W�2B��+��]�,�0h;����xf1 �d(=���3>�i�zwv�)�2������Շ@*�������}@�$2��w:�Vj�.`C	=gF5�i��քՔ�;�{�`%��gr5�"��(�YQ3�E_�x�!}����%��J��(�sAۇ8b��Ե;��x��ߍN/������]�c*+;����	�����4J_B���eԲ�9��yC]C_C�'k�V��E< 4&?zJ�Hj����%�ן�2�i�B��eV�?܇���Z��Ǿ[�5���]�+�6P�Tc�����ē[�v8y<�U���!�w�Z܊��6�V����O���ڀ�НL�D��ѭ�����1�M��	��y�����A�<_����zw����j\ܪ���*��Օu;��}�"�v�d�*��Z��_;�/��*?��j&|��F��>�9���Fag���?��Vm;)a�U�pR-&��<�\y�cX;}ɕ�h+�\Ex����B3���:%R��tGc){�����\��I���I-H���&�5E�6�$,�
�;��ͶS���Z^I�����I/�O����Zj;}g����M�Ζ>g��r������%��쪚�贴�HB��Y��;�ҹ���V����:i��GS��k��<����L������Z�J�5tsr�Pj��>H��k8>�O�]�`%?$�ZLjO�J�'��RP|x��
��wt:����쟈�vR�Q9�;N�<�lf%�<�-~���]���N��Tq@�b/�aa=1��'����@(�K�t2�L�6O�X����1��P"�2��M�{R��*"m���� ��ʏRS��_�~lW����OÝ�L��_�RT�{}6�8*���maΏu?�/�a�?-d�Qx�Ls�aWVQ	�rȬ~ɣ8�1g��mn�������n�������愦㏔�O]?Vܜ|�8JfT�n2�6|��_���)%��Q�QA�d�Lt|����	[�Y#}��+aB����2������u,%���G��S��SmÁ���)�P���8���)*��+?��vp�C�Q� ��c�@��ޠ}�(%��s���_жO]�Vpt�޷¡o8�ꌨ�HY��,4�u�0ߖs:�Sf��󯵀� �ƓoT��ƺ�?���t��{�f����ǚ�X�c�CO5W_fi��R���y��]`c�G��K�ѐ�nɞiű�)���*L����SSy�k���߃��Y���������"�� �]��cVa��=�"R�������)D���,�����u��i��  v�=h������k,o�ս�=�D�TL�QD����k����}�c��uXV[��>R_hŦ����_%���
��\dQ�q2Mp�����7���_F�O�C�g�E���]�H�v}V��;�l����{�^2���=9��[��i�g��J������lA���+��W�^`6n��^ �����N�Uu���-��Χ/�=z,;�����ﵐ��ź#�Y�8"��G�=KEO���?��A(�;��_��h�KG��8����ܛ�^�tO4�n2���z»K��2UjoЙUhZ�z%V��e��F�3~��#��o�jU��9�P���9F����3��=g%�҂M�[U$\Ǌ��=�����&k��B�!2g/�'d &��5Pf�h|g!��w�6i5��u�l�������+�))�o��O�x�([�d�ʺM��#z k~<T�f�����J���p~1ot�5��vp�I���?�;�?��<n@,�m#=2�RB�����3~���Ǒ�$v�����E�IK}�G_F�Ά��7/�<E���lf�����d�G��!F�s��$�iw�]���������L.\����z�Y)��k�p0q��,v���wn�c��`���XY/�N ��՛o�Ĭ�''�P*73����B�As1v#�es�,��k�T4Kؾ�����7�)`T���ǚ�$�(��t�xx3 �[�9�B�ϊ_�Ւ�y��s�����H���}�������a��2���FN�.<�`Ɲ=���	�g۷'���k"�>\�z�S;��?Λ�8ң��� C�8c��}آ
���+����*����^�*���J�a�3�)�w����{���[����5���Lh**|�N�e��M��Tђ�YM6�q�J��z�B4$�nBc�u�w6�M�C.d��z���K�"�cP8=<��y��X�5e��s���������m���������}��-
ک���L�Y0Y�&�c�-1���?x�}��#a,�|u%�m��e�<茟ͳM��u�C.�2u���ixkC�Ͽ�p��5l�w�U*��-�����k�բX?�}�x��O���%�:{8.0���P{wB���9!���$��w�5���Iر�����~'#S��y���Gc`]����� ���|��jŎ��$L?
�������(1=,?:�q���䴍�b��������{�<�_�Y�F��=l��W�y{)I@�����!=7��r�X�8^���?F�-�g�vn�_���nzvXO}��?��B �lG�S%%Q�1ozk�Y�ׂ4^	B��Z��3��P#�l����Y�L>�U�)�����?���;0
� *2�Fg__ U\ޮ}�����������EJ!΁�R`a��Ӓ������y���t���LXh}�}n�g�`�?�����-N�_[��r�T��II�2?{�h�@�k�k{��$��*_L��0hi���N�a1�F�hvH�?�3�ѯᖝ�����o~�zh�%���[p]I&��=/�3���ʡK��&qq=jl��)���)�*ζ��'��OL����3���lz���F��/�h}uJ����b�!�����Ɔ���w�y�Te�uB��~���a�o/C��Ц��Wn�p9�ɹZ�y.��H�Fd+�����h��y�.	���%v�����e��#�іMw�c�O����H���PUA78��@7U;��l�e���N0��������÷����{<1�&��y�� �M|�<�v�-
�z0�y�Um�� ��xw�����ė����u��e~�]���ɀ}��skQx���S4����_	���EU��4h`��,�k�0z�s�ҍ|���=+�}Ǯ��]����i�kc9B�s������ՠB� � �61"�v�\iT�I�-l_)3ߞb�!e���o��&��%>�(#�����ܫ�2TT����Q��x�E!)����^�On
�=$�0��M}3G�|�[�F��.��_P���{��w�i�s�B��l;�z-�8y4�?���-�P
���b�}5(�d�*n��=��7���t �N��������*Yx�����~��u�46��s ж��!�	�r�4�6m߿giu?�f7�	�!D�"g����ࢣ�=j�G���iGa�ΰ�h;T�Ni5F$��ɓ��j_��Q+]��1��f��PrKT�U�4}?�9z,/O%6��Q�g�7�:����][҉8��LKS�����&�hd˃�}}�����Ne�5)5�/|"xB�M1�T� l絤��L��������O}~�[-/7w�c%�WJYM��&(A�JuM���L�a5�6'W,]��H/��DX9�����F�x��������T�]�Ṗ�b��������,���}"7&�*�@&�	�4�k3��5J'���e�c���4���d�3�Ri��{���^�!�!!���4ϋ��Nv~� mc ��O�߶�O�EaS(ګC��Sl\��<x���>�d�u:���������B "K�����&�4:<ǳcsIO�Y,��.ͽ��A+�G�X�h� �To�\p�0:�=#ׄdLɖnb"��so�ud
�<U_K=
ҵ�%��~he�v�k%���r����uG'� d$���{]ZIl��/��duQ!Hc��k=Sn6u<������hV{��ek�V҇�;5뎀��KBx�b��o��1!�$>k��AZy@X�W��x�1�:EM����7@fq�[�*���}����d,�~��m�j��ez�e��g���{ތ�È��|��,�5�����׶���s0�0(�0 ��j�Z��;�3�λ:t���B/1�PH�2����;�{=�C&Z=�
����5"h���
�*���자��5�Ӱ�&BK��+��޶�%������W���<��H��'5m�Qri���� �����c"j��~��7ݕ��B�J/.w�}7�J��[�pڮ�D& 1�[~��v�tj�ٽ��H���`�:I�z
�y<����FG�_Gz׺&#/}��X�C�y ����s�V�P)�(�?9����%t���V�nDf�+�:�O�I�A���{y8_d�p��R����w�<����8W�	K�J��<0�hv	BG��]�;�P1�]Zw��-�X���q�IJ[.��~��Eڃ=ը��^is�l�=�^qpN��;d�F���usf��:D[ݗƽSRR������Akw��y�>�J�q0\P�>\�'xo�":AA���I�0�T~/����9wˡI}H�����@�w�-
4=�E��k�Ǵ3^�sr�����H�a�	A��1���^�%���χMe����\�͆�  \,7!X)!K���˂��L�C�-�&RR ���g�9<�Oo��fa<ʩǸ�Ϙ�%^�`o�|'c�ly���V+0�`}�t�+�`���tx5� K;�@� �
��q�-�V�y��儒[݌_������/C+�J<�}+.@��7�Lb�L.pL\w>�+V�FK�o8�5T�$�G�h���z~t�Z�^J�;����e��.yS�����W�M.���?O��8�O*Mc8�]DT|*Y��͚����}�`�
mmj�<{=b��QA���UI�o�nd.�3�M�^�����4c� bk1���-�q\R���q;��N-O�J8d�ğ�e�~�����;��ቀ��/����X���诈�kv&M�����\pZ���V]s�ŗ�����Q0BÔ5���kD�C�213gƧH��_��&�'i��x���\��/����7L��8|��j��5�A��
n9��a�X�ʿ����AE���f~�)���v{�5��[b���{Q$��x�T�5@<7�HG�ځ� 9�|�s�?h���s9�ϕ�<��k�y'�P���-��V��-���-~� �{��ܗP���x!�yS�	�@�[��X�m�c�uM$Z!x�i`�oZ�IY��U���Řv�O?2̤�t="��H���(�;�<�g�G�'<2ΪE���IPO������h:�N�ͮ>��Q����3�<��Qgr�a ������z����9�͙�vmXX,:���#*�.Qc9�~)�<-fx����� y�ϯV��nJ�m�NPk��nڑ&��G��b�E4�pa`G9'$��ǻ�d��Ϭ�D�08y�?2p�c�B�`����0��/�H8ko�"���U�����IЃ@$�M������ojOad��\����b8,��2����P���x��)!���#㵸ر�Q�X(��&�~'�rFΘYX�i�]����H�G)�r�'�������y�{��?F��|���#�9���i���N&��`�����8K�qT��E�hr��[�?Q.��!��Ȅ���R��VF��5�&��ja>��6���(��M�_ae�M��kU���?�rr��=]�Iُ�� ͘�A�yaO�}�Jz4/�*���b����I����=��ъ]�s�?�9FV$2�姍�lM���������O5DçOo�w��D+�Y�^*
O �s\�Cc�����E৾�$yS*����=+���@�R;s�o�c��+���SS-�h�<�(;�J��7X��ۤ,.{�e]*�k	�e=�$���Դ�"�_��ܫ��2y0m����|
~9�ޚZ�80��<�e�iq?���UY�f��8�oj�˰'�����-.W2n%�zeք] ���X_;�C{����7e���)��Ȁ�G5\��q������Q���k[�廜'O��_�	����jgCQe�q2�D@����ۭ+!kP
YN���d�ئ�}=�$��ؽrީ���n����?��Trc/������]F���ȴ!cw�lϭЏM�璳��4X�P��_e[�Ui�c�ql-�"Z���omw��������
�H�?F�xxI���P�U)��4C(���޲ys~����5�$ES�{`���"s��0+j��@�<!�'#p#��y_$��m��2���|o�~���ᙨ[�{3����q�ݥ��E�H��3����E����y'�i���y���WeЏ&�EeXm�
�~ӾS�I}Wy��`�I� �3���Y��[�O%g�0o�p�;��w�[Q��u����Q�xV�]���N�R|V�?3z�NVИIʜ�u�0���}�٩f0���	��hH�י���d��;��]���8��a�����ba-E ���\�?��m��������ȝSWo[�
��V�R1���<!��Pm��$kMPy�=q����	�|%?��5ғ''X�
[�5VX2�A��kk㼝��"�����q�$��^��@E��~�-m�ĥ�F͈����)C�Tq��Ü
:���g�&���!}]�,}�K�^{�`�9%{o�J~���Q�ˢN��+((2ؐk�q�;��u���_Z/zv�<��W��������'+{��1J���mw<��PaQ��>�%�� 0�4���F���Fv�ap7�.�f�JQ Z/�!�(�`=՜s�/,撲b��feH-3y���}�ɾ�5Ğ���(������=��
��d�"&'����6`U}r�Vy;g����PvƕM��oX&g��<�
ɷ����|u�\����	Ԫ��N����h�v�(�!�%J�q�94m���f��� �-My?$�/_\grd�vڇm	.��t; �4-7��4f�a֮�YIkR)0�D�|ҹΛ6^~�?�5����u���i�{QQ�:}2OFJ�fPG�[S�7��y�3��K��4�������K��)�]�چ�x���kKzG�K9LآP	�W_�ص����-,��K�w�&Z��u�*0�#��&��<é�Ap�D�>�*��O�%絓��d��|�RS�����u���̌��T�3�mS�������Y��T�0b�7�v��O�:�ޒ�E���/�qw���)��PE�:�ae�/W_@�q��+ف��b�&�?���`S�`mM��?����D�|���WѪl#5x�Y2�����ݿ�����/�����8��]uIO]߿q��˱��˺(E�\����q���-�\����O	&N;7H>�Z)�F��e��u�� M�i�]g�v1��H��z\��5:�U�����g�a�a;x8o�Ʒ�F�z�/O�(/�p*�[�ㄼd�}$Y��O�#�-�:�8*�/������k��i՚��)4n�y�����fГ���$Y��jl_}���Km�q���W�=��BA�����W|:�N�?,��Y�o
�V��V8Ђ�W�VT���a�c�+�_�I�.T�=�`(.Jl�#�/3�\/a���k]	��9- '��{�7 �pNaZ*s��_�E�&
#xyf|ZV�
^٬贚�4�4�u=G��ޡ�m�y���!lu�NX�4L/�b�N�˿-פ�ޛ�G���ܲf4j�uc��8^��)����9��>̧���`n~gVJ�W,8KN*��3!�� ��\Dlq��Nf�<;�kY)	_.�][�W{RO7�=A�j�'�qW��lu��eChՈij����'\>}��#��F�G����Q�SW����:4� �=	�a����g^�跾�қ�M'ĳ0�í��#���5������5�:�-Jo���{�EKi�J1(�S5��x��i�K����{�����S+M�6�]6L�ivky� [2҇�8�)�^^x�s<@�0�5��4�~mQh���k �{��}2�IZ4to'�`(RL�f�OW?m��T��9���Ir2c��T�������@vӯ?0WE]=����&S�yJԲ� ׿�����DY�»�2���:��uT�#���2��Jd��t�k��[=�K[���٤����W�P�%
!�:H=�e��v(�\��3H�,`G9�Y�v��X��1�y2����ӊ�w++�f�#��%�ޗ������Ё�̾Ul�
�c�6R�`����R�]U�Ш㸿[�$��H��5|ʌ�8�v
���*E�B��Ë�AcC�ή�Y%�B����\E�-]k�p�ŋ�Lb@�;��_z;;Vl����v��Oч�a]�����ݓ"�����P�h���l�;r��y\�Yû��V�7���v
S�ɽG�'�J,w�~�sј|m��}'�f�Y�vsm¤�`���m�'Y�gi�j(!F�|噏Әp.�Ojk$b�lU�=�r��u^k�E�M��Ξ��{�AaMݧ�����^�[3o��H۔.�������	||���Q�
�!g�"���Oב��&��U����s���-j�Lx7��_�ˈ�8w��Њh�g='�>4����q]�O��0r2����'Z@��#U��T���ӡBZ44:_�@�V�j�ܝQ#��-�g�Ⱦk���$qvC�dj�D(Ñ�Wa�-�MtH�uz
�uu��5��Z�HŖ��s�SmQ�~z>3Sc;�O��$�w57����`[T�#�	^�LoEyK�nߤw�:�bl|!̺�zdh(ϣ7��CG����k[��&LZ��,��u����߮L�y6�Ⱥ�����G>��O���K���l@����i_� �_;p��R`uj�Cq�����,���>��q(|õ��H�PK���O��ˆ|8\1�ܢ�t�sg.1c���:))�z�}���)�zԄ�����>�3<�-����]E�-��Lݷ�X.X��~4F�)	{���n�N�m2y��u�������\���~�����^����^�BT��Y(a�A��]B�(�#�C{�ș	������쭻o(jn�r�jE?&�Ř���1g7nY5:-��k�"� ezS�~+��
1��z\�E��Tݛ�qo�?���oPK����@fY�ǂ7X^��q��<��^���o�x:1r��Ꙇ��y�S��	�L��`����2q�I��� B�M&�<�����j�9�?�
��'g�{�(n#b�ױR� �?�R�ԓ�R�1�k5Gb��{���-�CZ~�����d�-���;�y���t���e�c��an���� 3IA�%6�:��}�g{K�H^2�	�Ͱ�yA�-�"�1<5Xdl�C���:+C��ؚp�:QFf���O�Z].���)q#$��L���9�W�w�K�Ͷ���ܞ>�K�ݭ��&Z���X& �[l����j��Y�ED�3c��--s�Nv�7ak����np� �Ce��y�w�Ma-��桮��/|�y�4�Ĺ��&.�m`�<��"~�f_����D{��˽������X�P��o�Vk��$薳��
T\��>*����YW��Fx�����Z�=�ɮW4h��U��D��UU�RfX�+z5�}B>�b���t(bfa΀�O	�Q%Ӌ��QD�,Ƿ\�C�uѤ'b3᭹R�3�Bp���$d�����;�Py��Z#=ւ��7	�XL�M��/�eO����^�x0#C����KiUp扊��<O��Ծ>#��N�?��~��*�J��C��<P突���Sb�>:�K�2ŮɸU�f��+%���X���M�g�Ըs�ԭL]���z��b�ReT.�l�)�B��K�^�c]���1���|8�h:	���.7E(� ���h��k�4{�v62w����o+w�����]�};�h��'jO>^jQF,�Tnd��ԛ�k4.f,��N�9���v�{k��R��l����qΒ������s^��vJ�X��.���Rϑ�����J�	�ح��`���qF��A�rO�L���K�v��.����>���dK/�g�����6�9�Ν���Z=��>zD��7y, %�( [-��p IA�J7�S��^�T;�M�%Z
VV?!Fzc.�������"�#�r�����SC'$&�8v����@�"�kM2�g����K� ��i�K�-�S�;p}�{T�TCG|���#<�|�9�5�X��8]'�Z���LyC\��D`�L�Dsa#���&��D�P�ޡ6����Y�Ov5s��X=��	���>ė���.:*(����hڞ��.P7i�\TOCs^�{ߒLߙ�
A")e���;�4��"�R�'��ͫ6�*���+�!RcM�/����G��Հ��]GK9��c&�d_Z�~�)�M$����W��kh���������Y��@��Y�Х�d#d �̶FH������ɋ�u�ݶ��Cy��Ek7V�L��9Ǵ�,�����s��6�Bk!�����/�LFN�>:np�h�3�4�n���;�|�o��d�$�
	�3�a�Wܪ*�����
U%� ~Һw|�=��`��P�O�??z���l9���1?̦�+V\|˪D�'��`a儁w�$sw��ʥ��&⏑Q��=Q��f=�*t���#��w9_6���'�4f�܆]}g$��3�>���j%'
���'�>�i���v���T)�!�d±["�}};�^���7��r���VV%���o�y%�c�T�+zRX�B�� Ua��{��_JX7�j�����L�.�s�Iq�=��sE��y]]xiQTXkԨ3Q-P�'�7s^˲�,��k"3���w�rg�F�B��6��S��n\&���	ȥ��9��"���2߀�d� f^�����7�O֏���&C[��;vm-a�ٲ�Z� n{����*�4!�UT�X��6�׹Go-���J�O>��"�`踶/\�N�S�<��=̗�N�"k�y�U��W�m�

�'�c����|�����߳��,��
��u���c��!e�JB���� ��
�$�#���9I��ǎd�=��,~!��d�M�}+J�o�u��x�߼�/#�������B�@��7��\�/�%d��+=�~�O,N��A��,�5�ϾtnGZ�"|u,���

5 ����RbiWK�<����9�LL��[�s+3��ĺ{d��h������Kr�@�Z%$��	c#1U� ����ڛ����H�.64G	Հ��%恡8Tjr����_�L��K�D��``�Un(0}��u��&K'�(��O��zl�z�ZW�,,��Q�+M��@�s��F8�l�����bgac#�]���ﻮ0�p
���-�r~�l��S�d�<�
)~=g�@����ڹ�^�ǺI�΍,�� �a��R&�=f�h'�6B��G%���9��W�Tʺ}.����ʩ8��WJ��Ui?c���R����k������:zބ��6������+[�x���	����f��o+ٺ�!� ���)�X�ZfU�s��(L^�S_ÿL|���ߤ���y����Y�3 I��.��c.7�Y����X)sx�=�[�W�\#���*e��[G�WF�ѻJ�{4*%����Կ���@�I8�Ak�a���z���w9���>zN!����J��,�h�*��ȸ��0\��_�ap%��9���.�.]���L��4|ۯ���܌>	G�J��ܚhA��w�Hes��r;���2l嵉8.�˖���R`�ڟ[#�?Ak��p`��x�Jv@�򽰳�}/�X�/�,UK���^�gb��B4I}�9�����@<����9���1֜��vu���m�p*3�V쑛��p�~%��or�e��Ii������?�����RJF�Z^/���*Vj���b;�6{��{�����W&�2�6���m�����/#�M���jo�n�ըr(�o��Z�vM����GUs9������**W�~
+��6�a*e�+��>_���2�}2v�����нﲩ;�	�+�������m��c���I�~_��=�^�82���}	�W�-%7>pӷ��]Z!�q�7�����cY��[�o�k����<<r2��'`���>��,���zf>[�A1�8�7��p�/���5V�M��3/�Ꭾ|�6�ӻ�=�
��$�
0E:c�U^���Z��ҙtt�TZ��L\_���,)H�*A��y�tw�?���qc����'*HF�L��7��l��z������.�>~�ssWV���>���<];f��z��n �	��J2��&��Jȗ�sX��V�a`O�V ��W���d��[�g�m��l�3ӫ%ƥ��7E���ԺF���&=�����\1|���lټ�AssuM��U�W�W�ޖ$�x�}�����|��O���8r�95��v��7�!&�T�V*�W�����bm�B�����DW��l�Tۺ��$�D�2�Hk1%����n�wOh��\:�L����-;��z�Ѻ�ݱw�����P�yM�=�C%�ٽ�a�Fd�z���7M�����E�[��� چ�}"?'Jk\��<����|���k_i���XiU&��W�v�>Rs~�����U�W�J�c/�W۱�P&^��g]4&���L��>4a�3�W��#���i��LT_�4���@`�n�:��*�kR
=L}<<�KȜ���=b��G�Ç@��Q�����XI�H;t�JӷU���������+>B��S�21$ZN95�с��=�+v��у���g4���o��!������G����"
�����eu�T��@h���bX���]&����
2g���F�� ţ!���V|�uC� n MeA��
Am*�E5�7N����ˢ̄���TIS-�w/ɯ�ǽ�p9���_�Q�
�8(��n���5��U9�Eg��ځQ:F�Yv]�������=�����	�>ܮq�>���#�A�#�e�w�_s?`��P8T&NN�f�����t���PF]9�<�ZY������C���z�M���H?�0���;E`��!P�� qd�ގ��P�ۇ���7$/��Y�-�v��_�G�o+K*Ӎ� �?����̮£�������a�5�l��̌�����#�^g��|D
�W��sA�R7����m]�@�ޖ�ں���6ΎS�̄Zpp�R�<q�ɦ0U3��p���P���-h&}�GN7=�c[�'5���e(����[h��=����=lӶԇ�����C�^���,�w-�q<�����������V�F����#����4�H��L�
���1�,��������vG����p�Y�c[8�2��nj�\�"鏲)(H���$�����(`�C��`[���{qЍY���vc}}W̍U<ѽ c�4(h���)����褳�2S��D�_A�8+�\w)��2��f����B�C�m����v� ���ckR�vR�b��J�!=z]�^�S���~/���rk�y��)�����|k�duU�UAi��6���u4����"��j��_���l���e��d�����ה��* ��	 kE4�\2����l'��o�#v"3�OF�@8R���T}��Τ����<�D���b�+��E�	�2���� �;���4O�n�o��r�GW,Mew�؃/Q<��ۡeW)�x���]��߿���Q����7N"7	�qC��y������|Ie"�ץ8Tp�豭 1�*%pQM'd��]�´(�	>L����G�g��S�Gө�!a�+� 5��/�n��/A@�vb}�J���o+��hV�����wy��n�;q���m�i^ߓۼ�ϵ��L������Ym��,��tTOي��:|s܃��z�(���6�5G8��'���"��dB��=���uj[��@o-�$���͑l;>"1>ڠê"�`c$zљ�L�y��䷎�<���6F6ٻ!D����FX���O���؆�� ��s/��M�?n]<42^�Wtc�(���Y���FP$U��`�;��c��\:��	�l��w����ݒ��TH������B�g6�����iΣ=y�<�LA�E�L/�-L��ib)�ٝ���^8l��B@b���uE �og�'���������϶Oe>zP�>|ؕ)��sQ��,0��:�.��y��
�
����:��წ���)��=�&�A���V��G���>���?��O�>L(����d~J`5��8�Q&�yߏ��ŉ�'����Vi2��q�(��Y�Bt�W�?���.'��d����(��j�k�;d�-Gbvefs��qd����}�D75lˡ��-@��>J^l����`�_���a';�!�wW��F��M�ۄ�K�u	��Kc\���ݚG�Jim^��]�V�Q��.��g�H�>��;cy, O�Ӥk�E�v���L��K�OpuSnC�0��Є�����E_h���síl�o�t�|�p�����ƪ�=�bb�����c-[����N��bR�u6��y��;-�[�S���~v[B
I��y鍔[E��{�uh�^�@��#˷����[������,��RʧA��x�lj}@��5�ˉ�)�J�+3�R�X2��6u��}��W�P3⍢D�#���'�����@�2�6���=Ǖ�&_�ɘ`_��9����L�{�U%���q�@��-e��K����ns�#�e�ھK������!������\��"��1�9A�����0��:�Ӯ�iL���ŮYJ��$eL�����q���Q< I�Ô�1��QՀ�>�q(��q�}r�&$�P[�C
ڮ�O�~�Ů�E���n�"�!#��Y}�}rE��:���e�[��N�����G0�.~�� S�%VΧ�j��\��&����3u+��'�-��k���'�`�[	:��/ס��b��f3-] S�6Λ=)҆*�jX�D:[�~k�4Inh���Qioi0���_�y>P�z��Pp�Y�������7�~HQ؉s�3���}}(��x�M�?p,Pk�;�/�R��F|*(���>ej4�����\n��ԇU�&�6�%V�y�I��DW������맪f8������U�ep�IK��7�.�����+Wʨ���C�	o4�1y�W�OG˂��,����<b7v�2�o����I��?�B���Ne���-���X�T�r�qВ��W�q��+p��BF&9����5��EE,�y� �փ�9��|ĺw��K�o��G�*`ay����m�+C-K�����s���aՎ9����z��ss�O���� 8�fՍ��I~�4��W��Aގ-[HXxlK����_�
�4P�'Ykl'����Y���yS��E���b2���UԷ5(Z�q��e:��m��J�	�����D�:�{���}_ǌ�og��^� ;k]��^��$5T��t��ƄH�!�9$�5�e���ۥ���
�WN:Q���-��ۄW�K���29.�������ǖ;8��U�
"����������sq�������d��;:�#�����+H�&�A�j=X�MzWBG@z��@�%��z�gF<�������r1��^k��^�}���7���X9�HK�+�ۃ��;u^?�s5��p�S R�h�mGX9h�m�rn�����J�=I4�Bs9L����w8*X��'|�5::�����%����%�I�j� v�oP����M�`	�e	@(a3X�)*Z&n}�ɉ���:A�,.W�����R]/����ğ'ih��]���qr��|�|�Y�ڎ3��&���p5�`���m�f��4@A_)��(.��,d�ѮNpȝ�3~o�pF���vǇ��7�~D~���9�������F0�(4f�ٌ��i�'��_�@u~��yI��\�xĉ���{ ����8
p�s �\�7��|���㼊�Q�'j��N�9�&L��{�o"���H"}�Y�x�e��@�	v�*w?����P>�W�O���绶��#=�l�1�3������>��F��Q�$^��}�'l�ǭ�׃�cm<��P0���s��O!O8�x�'*���F������C�s�X���
Dv��@�Ni<کP �>(�3�S�� ��ZX���=4�o>��fb-mݚ
��[� �~̽����
�$` ����ª����g����f�|��,�/-KCw�o*z�8�H��+'��[K�5��:"�3O��_8��S�	��� T��ym�B��� �À��᪺���r{�3,���t���ֿI�O��T`e�YN���Z[N\E��;����N�o�8��{7�ir�-��x�i��]	Y�bŝ�Xҧp=����9��4�\��x&�r���6���Q�H� j�`b'��G�%����D5Ի��_W��v t�)N�'l"����?߶6>����� �/�0��z�Щ��so�F}k��+�}%�oON(���tv�t��
�6��-W��I�����|�[��Ք���Oe��#���N�<�jL��~��]��g�D�a�����:�|]�-��$O�-�p�t����Jώ-��asNr������9as(]�z!GOF�`�G��9	C���%�9�~���\J�^B�fߚLze�*S�i|݇���5]:忳8�\=� ������n��p���#� &�k�~#�IR�s�6���w�U�5b�PvN��.���o^�	�7�ȅ^�����i��_��{��9�*�zz�V�����ߖV��UI�<B�:�Y�f!˵�*�aXqX�_OK�iv�8�+>>A\4@;⻋����&��ZCX��'�|����e_翿9ʱ����x�hzJ��D�y�m>l}��D��VD �	CE���MsN���h��{ߠ�*Pt>�jK2|�qL��
�SQrYE�d1�Ψ��xm}W_z3�So��
�Q�[xY�x�S�"_��݋����q��B֕�r�2��ċ޿�ɡ�X�f�x�tF����S�]Z
�yз�ϯͿ��P){��qj3����N��$���o� �Q��ZE#�D7�>���O{��ԧTDvܳ='��=�_%+V�g4�i�s��o��W���Wj�z�)}�|]�3�j�'N����ͨ)�סrЗto��|��r]��繹���kri�!m2�K�2�6h�����#(����Ni�NM*v���,低��^ f(�l��J]����E���f�q6�\R�p������u]�7DO� �N)(�8��s_��*��G��M��<����wD�V�����.g��������G6�0���
`�m�rC���������:T��F�:_i}U�-\!TޖTa�׆T����s�h��338�aE�(��7u�y�`Qx��MV!;�s��^�pvrť|>�%��W#
j��}i}�t,�qJ���p�t�\���d�4��)썢TrK��-x*y��|֔�[CCV�D�ia�w���͒;F:��0��5�2z��%/Z�]?�xR��ÿ���Ϲ����pO֞�HSdm�W@e;��RjʻJ��"�/�~����5M�R"����P���;�9�竺��V�>�w�q���lb^j��c��w�SS�������UNK��N�����̒����#''�f6������2m�R��Շ;��+����(���=R ��]]��E��������i5Cx��t������ތ 
s����|%��!��4�f�=S@��ُ��W�+\l�=��u��K4�he=j#6x��sNSƚ�.V������pF�Ԫ��L:�z.�!��B��Z 6��	����K]��B�b��nG�]v�4� �/gd�j�(QO�eiܴ�-��eB�p/݉	|�{U�)�G�+�XC�X6�]D����qmc6O����{)^M>�'�ϧ�B:�n��/4�\vl[iu [ǥޤZ�\��9\�)Q��EaU����8���b��t��,f���3��.���>��[��L�z6����饺�_�9sP�$��B{+)n��ԗN���y���S{�i+z��*�*
P)N�V��=ܒc	��ܛ���*י-R�u~}�bhY��D+{�g� �YP1����{+g��-$��_w�)�*�%)d] *5��J7��f��v���J�^��׏y��y�;RP�gm��$�����x���TT�V~+��⧸�Kg���}]���60x��i/{s�pAj�����Xj�N�ՋʹNM~kJY6���#�6e#m�i;�sz=�H�l������T�.�<?�YR8C���>�I(>A��h�L�{����[Gn��-�"�W)��kUJ�����:O@Tު�_5
�&F���yiP��,�%��.R���3����#O"�bqn��9ǥ�����J�A �ss󪥛��Ń>�|	�g�e�s��y���\;�Lt/7�9�}n#���f~����/9kFz��g���θ�����k鎗����k����L',�����|��T~���biq�J��ܜ0�����,�n�	|~���)�Ţ����VIf%4K�en�Po3j]��*�m�(s:�p�nP���r�~s���k۴j��{E�f��=��jhkS��4#D�4�]�s�%ר���Yn�� <�D��t������鞙+<� g-)���
}�K���'_�Zl��&��3���U���s�����z���̉�HË��k��#_@�~�����pk�)m����֋�ͣ��	�J3�<{��M{��E�a6��k��l�����wB�pw�L�z��Pd�s~g0-6Br>�R�5�#7��HӻeT�c\Tr+�,#�8ZW(UZ��ܸ]���;�_���(N����ǁ�>��R83�g�n8X�L��Ur��7v3�����F�f�!
�ˋ��p�j����[iw���{Ro��FgqhoE nҲ�F�s��u�l���(gI�d�^1�^G����4-�p��e���4dן�xYVc'6oո]q�<�#��痐���/��������JJhԶ]a�)�Ǐ/�a�قu;��l�T#?��\��&���pJ疕B��ޠ/�ঞ��k#�/}�J�K�5��⭵���L���cm�Ѻ���i`*_ܼ�u:V�a0�Ǘ�Dmn�����'�%�٧fN�7�2�[��5�O��"�t<~���*o���r��C������1���9=�8�����G�h������h~%�ǳ��-��O �p��b�����w�7{�~�;r��?zH�C)�����&�)|����B\��˚t>�E�<:6�l�!+�����/:�p9T�t�����v�R�P��.���XA}TQ���!����R�9�X�_��.Ç;��^b��0�|�ȭa��嬎���&>���7��W��{k=.��ig�jxu��>0�1�%Ct�y|�k���D�F�bd�p#����q�q�=��2&���,F�j.�=J��#��ֵ���L�z�1k�s�7�]ʃa'��0x��5�E����HJJ����4�7<[w�S9��.�{����
�Z֯���s�d=8�~��Ul�sNr�*��TB^{��y~+��v��6TATFn�����#��؉6>4�FZX���Ъ�_�6NUrXX�뢫�k����<x`=�7t�0�Q��88x�z�ͱ'c�{��͓���_��o�i�ޱ԰�G��w-���
s�p�ZOʔ��8�*l�Wy%���?�a��|�؃�E���
d�{�1���9�1���Q�����d|�+��Z9��w�>�nU�"�ty�DG�&Fȧ��5�|]�[#�>����t��P�ܗ���fHf�.�~�2�)�$��!�N��sF�~��X�έ����l�$	��K1���yx������Uʲ��͑v�}�.;��}����i�����_��si �Z�';�������n�%�\b&��f[���7a~�ܵ9���\O��2Z��J�1��'�ճ� ���8��眺��\�KBw'�?b���(>�-F��F@-�����0'|2lH��?[�d�(JN�uP���U���j�]��3��2,�V*_ʟ�u{	j�D��&`]��*�f{D�pKD)�P�o�2�C��w��/��ϴ�j ��%��.8@\¡"��K}���M��CS�/��U֥2�
$����v|�̵=���pw!Kt/����c��Y����U�Fȉ�Z�.��&aM�+2���͆���zit�_c�z 0S0I����kjGQ��_�^qY�ǚ_�V�陏�-�r����
k@/�2�=�w�e����\rsͪ'�pp��R�_���^�]���Ww�u󌷧�<G�ڴs�(�c�xk#"y��zȤ�ɳ��M��p��g0��v�ho?b�������@%�$>͟ي��Oh�7�F�%����ST4�t׭�e8���L��m&ls3�_�h������#���>JW�!@���|5�Gq1v�
$ไ�0qq:���=-��j�\8>K1 |����ٮ҂�C`^�bbN��ņ3-}�K-)u�v��=B��//��
�][i=S��Ao��s�%TFn
��81�;?��u��q�b�|�^K_�vh��L���f�������o�Q�[XS��7�C}�U��tS#JI,�aW	m�@�
��R������@�m(Sv�=�ytx?��7���kZ�c�띯K��뢡c�_�#zAYV2���u��P��ڳBf��IC �[���1���c��RG9|\[��$e q���B9*�5{j��0h��f��9HQ;25an��"맛�w�+�؂��e��ݍ�B�r'm�i�3�=��*��Waq��Cڈ�W�Y�<�zur�;c2�v�e�#76�剗,11 ���fOR��\��%+���_��Xz�����i�I���Hx����x�����z�{ҫ�	��zJa����T�w��Q6=�������
��:��n���|Մd�9�[g�KKj�*���>��X�b<כûeN,��L�*.�6-y�������J�r�ُ,���� +o��k6�5�:��1��*����z{�l2�2�\��9OHR��E��c��A��Y�s{�<Þ��1���c�N$��/��g��^[���Hd���1��{�͗��1�_��O��l�E��{�#d:1pQ��W�S=5C���1Ŏ��'��wh��H�K��{,��JY���G6F).Y���*���4�&2F�?�Fc�$Y����S��h'\�����
��ok�+��\��������6�m�y�i�,��Ph�[Ë��8d�Lڮ�R�h�i��"O� d
SOi_`s�u��oY �]h��7����*�
K�[v�9t������C\\��1�Z߄�Ϗ�\|�ґ�P<>����Pv����U_]�/�[0oO�U*�]�Ž�=�86�+��[�.W���r�Ŀ=������#qo
T�����)E���NҘ�tp
�n�d�=��4/����8��B�9:����7��C�#=�bD�9�	�R���ph��ۣۚ"���fչ��>X_�ă����_���J���ŭ�
�Ш���Eec�|�v��Y6_���R��+���p~��$GO�Ͳ�ۋ��z�%pߗ��ͱ�F�ӿ��;��_oC��<v�rM_�7�Ȳ��g���m���-R�;zv�����-h��� .8*��	���q�|K����
#g�y��2n%�I@ ��^����9_��e[|�Q�`�RSNw�r�A��Jca�͟�퇬��������J9�LKys1�`��➕�6�CC꧱"��r��ND�23���〽랧*3L ��Q���mng;��7P�u��բҴv�7^@,k��/�ܧQ(��d,���{3�a;NR0�r0�u��c��=U�-����h�Z..���ZqF(ZA���ʺr���E�/Ĥ�� ��{o���z$yѣ⛗�-d> H��.*��~��S�E��5���1�^��{M<�=y�*���<S�XXN?i��R�#�R������C]^��!����9�����g�o#�����-OOym��]}�6:-盰�����|h���o�Vm,�;����������`�qEZ�U_�������	����k�����z�}\E9פM���5e7p*����]/�2O��GuzQ,Q\͇i��0�����k���m���6�@���K�)�*����\j���u����w^�y#m-B��䔢y䲆~����A~���	��)�Lsu:�!��:c�I|}S�.~9s��v<Ztwe�a��mc�ڥQU3��B�$]:��m�dtM�ao��S��������D���b�A�"
�^GJ���Ui4<����(b�4�@_�af����A)�,���r2����ae}�:�Waa�@�qlBIpj7��6z$h�./'p���=���{��&35#f��Z(9{��b=G-��CG��<B�b�u���$�u�gC����[�lJe �*�2[fY�g��\���J�eO\�G!>�aѦ���-���=_�d_���f��N����u�����$�Ϟ�1�.6+�-&����ftK�����iI��\U^��S�A�ث�ùy�T����i
}V��ľȿ�n'�C��Pdi��V�sͲ�޸Bj
���\tM�*e�2P��Q9/�[�ͭ��:^Gov�N�C�7~���mA��ъ��7�o���%yD~���A8��q�3��μr�nn8��v�9���'������	�<�(�X�̊��+�WJ���=}
����y��q���Y�����_%sp�X��R���E����I?�Q�s�`������]��A��wJ��R��a/�+N�4{;F|�m������d��W)m������ǣ��f�c&GN������DQ�PXVV�ᬁjUn����?;��}����f���õ���5yxڤ�LS���n�HP�t�;�?�tB��1%�vEݼ�T�l���W�5r�O�1�t2�Z�ܼ�6�������pi`�Rx����x�ľ�o�?O*I�"��x���8�q�gynu���j�>cL]����gyyy5��ϟ�w�g����rϬ�w��/��ln[��U~�� Ť����v�}�u��^��"�YW�U��)�s �%�j����D6�l�'XTn5��@l��/?�;�-����Y�%��V�s�o?ؔ`kj}���?3E0��it^�f}�E�F�����gO��A���?^>�j�j�k�+.�w�FTߐ�����\k:��Sk����w��(9 �iB	$��Vk������x��V��Wc�u�T�U*�M9���YI��j_�l.���8��ʂ���\������f߱�$�9���9�ǌ=��
jȭ�wi��O��8��|�@Ϛ��P[%@�S�R��rK��|w�e��ć2�WP�!pd����bL�\1������:�k8�#QoL���s�H���TJ���Y������PB#X�;�wa��Qyu��pLai-��<55�$dz�I%._���	LF˔��u�Bl(C	���sV��rN��F�r I���-�p�OI+y3�.^��ǧ���;��Ԥ��j�)�����^����Hަk��Z�����f�q6����}%�3B�-�N���0]�lHH���N����T�f�����܇8l�!MpȲ'�r�mZ(z�U���WN��m)��I��ԍ�y��)�gа���[Ǜ1���%"�q��6&�oψa��R�Q���B���<�L.V��O�׷y+���{]�vH�~O�%��!����e��7�1�n|�[7�B/�j^�f&%i�L)���,?�q�l6i�ⅴIH�csꉯ\��2�C0Rg�l y�XT��l>>�/�&ƍ*;uJbogN�������^
f�+4_~��DNj��V���:�0�t�y�}�/�5Iܺ_+�s�~�ɶ�;���έ՜������M�w��d��gҍ���MY;�wj�~J��7c�&��O�R�60�=�E��2��Ÿ�+�~y��# р+ڑ{��h�O� "����k�ۨ��!S�����_sD�gw�r��B��ؼ��WJ�S�G������ޒ!�hc�2;J���>���x�w����g!�����]��H�Nmd�`P	��Nf ��z-)l�q�g 4 ����"�t�J�����?�>T�Q�`b�����r�5�����R�cS_��TTI7|��d���X\0ۑCҙ����p� ����O"�6wT`��v�;�E�8˨��z�;�[�zI&��lI�Q��[�[��:}i��� �ӶWq�I�k{ύg���?�u+8#@�(�� �B.b����VS0PW+5�Ch����J$�ĤFH��pv1���Z�\16!U�?¡"����o�~�������w���{��j�KYJ��ZO�Mut�������?|>'᫰P�B��4�녫��wUǯ-���v�k�0�xye�0�@�����O���~h6�6.'K���w��x#��p�a�Jfw�g��ň o��^�b׮���=�~��yA� ���M�������Е���9�ǃ��ۄ�q�a ���M��yn/"�؞�tD}�ɳ��n2��TX奠���ϿD�����L�-0� ��}��'���~0�1�q����j��_=`�$�`�~A޽��C����߯���������������z0�I.|�i�)�JA��`6��|_���M��J�ȝf͟�6��l?w��c��<�h;���{0�Ն�3p��2���
Jf�ӝ���?�ʬ��$gV�N����p�P�ȍy�c�-��x�u=���݋�S�7<<�g�C�7f�����܃r��L	;>(2�<�e��d��y9��k�8l�D�|���Ls9�a��O$��� wG�>����	#��P���6
 mbC��s�>H��t�v�^AVb���,OA9x�����[���ܰ�MQ��%�C
�?G���z�-;;���o�{����J�@��JG�iq��O���W� ���� ��s�Z���q-�Iޤɟ4�Ώ:���'�� )OM�Dό�;���-]�+��Q�M��0Un��o�P.�P�� �����������ab�Ә�����M�81��z�]��2�2��l�{t[�#
����\_�O�_WVV����)2����Gqƻ3<)"8o6�bĿ������O�rD��*}�aD�9z��(�|n�"iL�jfc��IQGG�8#"3J=�K���٧I����nɂ�����uN.��{����0:e�����
��a�Ua)v(//f�Ġ��!�3�W��-Yi�x�بhD�4���^M]r�b�� �}�A�����%v�e��2$ޛ��N�I`����*B��_�^o��~nY4~��k���7�2��ʉTډ1y���y����a��q1C5T�ݘW��˳7N�(/#�'}�..%E�H^�}:��l�y��,��t�]W2��Z8w�TW�+����y	�j������jN~���,�-��P�]��Z��s������i��W��%��o��L��Z���󀀍����i	�9s[� Yu�^�5y���w[j�=�,J.o��+х{х�6��������[��դN�!��4�\��S-=���4����ܠȄg�����[)<�NYcn�Yo�IR��HH@ �۪�3�;�^���P�:��9f%V1�z���L�R^�%���\��(���PA�D(.n�ʙ�'0N��z�?��՗'����@#���;D����꼽�a@�4��юo�q��Aԡvfr��5d��LS)�B�:I�{��/��o72u��Ȑ�<�)N����p�	D{�/&��ag�i%�B���60��g䎐�Խ����!�Ơ-�%xE�W��� �����ug�G�Vr�K�n�{4��.ne�5S+dkD�"fo�z��$;N:a�P
�Q68�8S�QȰ�^jԏ&v}N���V��VHe�� fB �E�q���ӣ�D��\~}?�S���!~��l>.򸦣� ��z�q�e��_'<SY��oL]����_����ĳh�ʫ윜�V߂+9���w�����ws�O<u��\L��3_��P������vIJ� ����}���o��(��/�Ԥ
T^ı�޿L�\�@��!�=�D�Q���Z�{�h�����G�쯝�R}�bN�{g��������-o�}磓q>s�Jg��?^se{�[�$�M�*W��"���Z[W+��Z,5B(<9����,��h���(����n�*9��5u��;]g���cE�:fH%���C>F���X���>V��~��޷˳
���BL��{;i"IC����e�E��G�e�A���OQ�,*�V1�h_3�@�ی���z�'݇�#&�i�,� �{T����E]9�0c箾��'1�I���8���;���^K��/�U[�6�)_�.|��z�b��I����p���eO����\	2F,pM//Y(����OX���Sxkp�@+A9���08Ed�`|^טC�� ���>97;;��3D�-�BdJE��5�n�~��?x-e_T�cr>�չF���Ut�z2�ޕ��7��Z�fte𗋱������L��Ɯ��,�#.7�򢒐ƕ�I	����&D��6iW�3d[�E�P�I�Q�=ʽy"i}�P�1�<d�}�f���5a���W5`I�Y�̛Mm%���}��Sw�S|1ߟ��5�O��<�頩Zr�M:�o� ���j�+^��o�u���v�����0uߑC���0�>��C�ζp!�"x��ܟz-����_��/mxüㆆE<�3�������b
��Sto�8h���ˋ� �\��'��K����<������rS��U��	�,u� �I_�t�0�mWOv�~���4EKm�/F�%>y�ٸl	?���W��.�,�y�M�ջ�^�TЉ#�ڵ6�LÂ{���]Lֽ+&}�nJ��K��n�=�h>�a��L��/��f��f�Fh}>�_�G�5X�#��� ��N`�������{Z������$���9L�q�2qM�dy���S_��3��s���l/_N'O���u~H_��ī+����c�?y�m����M�����&����@V���������������+	@^!�lCS��K82s�r���+���κ���3�b���2����Y#9Rs����T�^]���9M���Ⱥ��g�������>6����g��#�CG]���)k+.�����v҂2K��ܖm�MWH	��ɸ(�Ғ�5n�7�HU��A���4���aB�.|�P��O���F����/-��抱1;j�,w��<�93�_�wurGWn"����7��lr�+�RA®���ß������5�1�Z0���3ty��|6�g����T���_RJE�a��z~7dN
��m�*�@=��u}�ꇩ�{�11�rn�&9چF�{�-����b�K����$|����hOg#_��rD�;F|sM�YA��	���g����餤�}�tS���x��Ӌ�����3dH�^�8Ѵ��_�j�N!MNL��a ���K�o_=W�Æo�]��n� ��)'l�hi�����I���P��X�AF٪a�Z���d\[K2�ߝ�+�2���S��]�[tU��}L|ds�I��Æ ߡZL�Ժ?Gr��BD�w,��.o%:L��,�����ƿ�b��7��|0�uP��A/���y�ds���J��=��a�=�K�`��L�U�	X&L�h\����L��K>n!���"(���@G��]Î\�Zzwm�f�& X%1�q�.�<*U�̓mt^f�Xb��ykl�rYVFa�����?t{0�ơ%���ˊI�뺠>���k��d�E��6;t�)f'~���W��m�'L��1+|!�ah*��B?�U��0�s<�"�����t�B��5Y��+A�v�5�v(k��f�a�6f�vsm/ōM��<Y8��#�׷ΑE�ڕ+)�`�ۚ0�E��8�+�g���Zx�җ��2X'���[�}8�1Y��Ӵ��wj��UTS��;Ni7���˗�5ٕ�e��e���]�6�1�:��9H#�
�M��k�m�r_&��#�M�;�����cw��h�+#s+�M�^��}@�${�O������'T	��I��CS���dXDK�e��ݮJ��~���d����	�+��?��Le2x����������9���+X�D�z�(���y�Nrw�;���������}lu���� rݽ��b��M�#�dc�L��1:���佹@�7�C��8Z�hw���3K=Aw�o��=�V�����-�C�O7��
 &R�6�������	�-���Q��2�F΍�l��=����u�y��&�����8�)���9��ir�.@��˸)zS�����@�>-w��r��;׆%]�eگ�L�/��y��MD��~����z���8f[�4�L�@=��8���:>kN�;Ϣ�k�3Y�cX���g�����7���R������]nQ���uS�C#=��s����ϼ�Ƚ13��@� ҘJ��J�!�o"Us_NI��}��o��U� b����:cN2�`�Sɒ�X �!��5K�s]��F�8iR�^�-����p�N��g$(D#��X@�O�wT~�ԉ�b�&��d�PDF8{�!މ�X������1�B�,8i����5�\Į,*����V�l6J.t5��<�j����)ki��%����,̆�U{�O��t���V�ߞ�v�+?l��ˀh��]LT+��:��/ܽ��ꗝ0E#.	��T/�a޾Pa>׽V�= !��T?z�8�!�1�ӏ�23+Z���o-ɉ	?x�qN�5�N�\�Ї~���lWF�1�w�á���=Ɩ�J!aG���&�;fJ!sy�F��ŀ�h��
F�I33���J��*����\."Ϧ��vw�t̑����c9���/�R���/�LY�����B��Ҹi��(�r���imUOBh���Kr񥾂��I��
C��f�vK�
�� K��&�~���Q>:�G��m��|�`�LF��nmH�0@C��c�f�cXIϒq111��콑������f�"F��-��P���]�w����X#u��VT�1uLZj��6�+�ů^��<kXn1X�+o���,Z�~��V�y����G�!l��^�W�ab-�L�t���z�����ڴE���snD�#��{x�ʝ�w$t9`i��s��=jѪP�f�^$R;�0���9h�\�R ���>�0�1�T�P1_�k]�5��~h4�����j��k�T#�1i4 @��}�c>H��\��G���x=�j
XA�*��h7!wg�j���ߪ�0�7�cK/C��=���lo�r��d+�2�? ��.�U��_:l��se�-=�0-y��������uݒ��)�I�rI-�.Vh6	��=�BRd3c��&�^�\���_��FR�9Í��'EZP]�����k�{n״K-u����5k#�6��u���Lԏ%%6���k���PGġU���d�3��P���㡪�7�N�A�D�*�J/�oK��7��!\�~
����TX�[w��j��`p�Do�t?�FC��z��/+�w�U�^��)\;��8΃��'�B�k�����	�z_�݋�b�9F�!>���CU_+X��}0l��D �>ZI( Ako��N���s2o��̋�ϣ争I�k�'��f�o=<����ņ��]<�!��7.ˡ�pY�
�!0�Vt#	Õ�D*��(1��L�f��Zs���`^���6�liD�v�*[4��[�J���#�u�S�h\O�w�m���uZח�%=|Ay�m�ث	�&>�ߝ�;+��̣w��}E�e���eJ ����ӂ�o�}v���}A;4n�~�IU>S��#��	6�9ݡzGQ�x�#U��'&�HN��|o�2�>ޥK����+oLq#�
�*F��kf˩�!�jMu��jk�F�b��^K�(��W(��
�2_�;3?�X�SY}�4#_V����4D|X]����5��09s�4oh�NL	K����㚦ebe�s��_T2mj�>��/��Gt�۞�-,��0Z3�d�ξԃ�`j�(��̥����~�X����w2�_r@ϛVM�=��m�؝�=���a7�p=�"n5^���NSS<�q*���Y�ﮥR+��$S�fDdƱ&�4٫3pd���/���
��h�t���REu���K)�~ڙ���(B~:�K�xv���~v깚�[�}���J��h��MDP������)�+ŏ=f�������!�(nT��{ #�yé�*��Ċ��E;� M4͏U[b=-��d���L��Й?5�
��9��L��.ϋ�zjc�،?h?�ͺ�*���|��^�.#�ۂ��j��"�((v2�,���9�!�ē�x�����ga��ƹҙ�d���KMıq�#�%W@-��gzK��F����$|�!}Z��ι��q ��/~�0�,�O%��{�d"V�w���֓*U~9�5p٤�l���i5��y��FW�ՀW^��A}���jj�+3m��:����D�v�!�.��`���C��"C��E�S���-�c����T.�&��qLM�>O�H_�<,{e�d�}�t��K�z����<�{9f<�iq��lTu'D;���� �b=�agT��$N��Q���ˏ3�N�U��,i2�d��J�v�C--����������oڏ�G����8Q)��\e(ki@�8��=t���AFL�R�*��(��H�3Buo'G�*������z����*dΨ�|��U$��{�!x/��f��$`y8��V�F�׹��˷�#w�R���(JcpX��O�����t��e�n�<~�nb�\@�,��e�.�c@�iLW����>Z5�1NHV�ps�gPf�ї����w��5x�\"����b��ZE<�ů&K!�J��8��v������^��L�)�Y�o�cy*�E�g��?F?g�Z�U[Cf�Y@>�쥠 @��m�4R7k������	&�O��_`�]r6I�Sֈ�_�<�!-����~��~Hvk��ͦ�c)�=Oמ�nz��P�,R54�?��IXPI�I�vX�"��V����ee2y���h������R.���������M/Ue�ݵ+6藍!v*R�ƀ��%b5e���ő&���/����Øڛ{B�uϞ4ZQw����<�p�}Ȯ4��}��5v�E�����|DlN�JՐ��� ��1\a�ӽy��b���N�7Y��Z���~�Ϛ%����k�'���	�;~|(��O7�w��`�\�N}�OY���h)9w?*��TWM�eO�XŴܒY-}v�ܖt]K}�8JY�v���I
���ZQ߂�Lk޴�ς9�Ƿ)k���̩�HT(�������[M);�.����3IX����8�Y�u�\r����|1@�'�c
ab1K��i�N�� �2��j���LM���h�wS�o{�۴�d9���(�}�h��l��o�j/0�Nh�7e��נ�E̾�ҀdWB�JC= ��Ê/����T����d�#�-f�A�z�8�
՚���ʞ��m�(72��!,���O%i��̥G`���/���9n����%�?B�|��6z��v�z�]8�yq'��v�.� 8�/�I�J�������AJ�T==a�۶lM�xF?���.��!5&�-�k��3����WaJ٤��yfd�Q78�����{-����.��[�z�!�v6�+o5����p��y��枺M�:~�
�3��0�K��K���Uߥ!�Sŵά��oJb10w�Q�b0�
oS�>>�J'�^�<�+f��3���UhXA�~��'BLC�(6��l��Z#3� �*�5�����:�!#��Q����lMd����?xgC�h��:u>i����k�fb��Ћ�Q�����s��W��fӫ�CS�s�����[z����8��8E���%������پN���#^M~7��6��o�?3oP�ۅB�����`׽&V6�����?Z�=�����#`���ϴVt�����SPX�x��ܤ)_����ʬEZ���7eŉa��b�tB��kߏ8B��
��tϝ��?�y<e��T$h6�{]�mi�
���X�Q!�J�[�w��9���A�M�!�,��R#��I��z��Y�{�]`�VN@�P�xv�Tc����yA���Փ��W��;�'���[�%NX��@�IrM���5�}kӁqjp�s��xNfl�7&f�oi�4���M|�Eǩ!օ���,f��1��%=L)&8�Yl�x��5a�����t���!��w�ɓ��@��?龻{��RI�����jÂ��U���{-���Ú"-r��J�5����@ɶ��<�^'W�e)F6i#{�s���#sk�}bǩ4�4����f�c��.�su-�'��݄y���&~$Fӏ	Atu��6��m(�d˙�^V(�j��ؑ�zE�����٠�BD��=�G�����4.���oa��-tI�=|B���3c�yM\�jy@x^,�����$Q���ЀG���R��Û6x<k=��}�䆧ԣ�.�~N=��.Q��]-d�+z	���if4�{W�/x~H V"ˬ��
ic�����K��/�� �;�qq�TTr���
	��Z\�@~3����hk��ok�U�JsCE%���OEq��u�j�ܹ��E�����Gp���O�LD���D �L��}�r9��w����O�g���~���(��%")�~�>~��s;�8l*�%��ЧYYg�ʎ�����uq�0p�� 54��,�q��>۽M��2�Kko������:.�y��iiii���Z��AQA�n�.i�XBEZ�إ���Yj�������?��]��3g��5ל��گ�2z��si<\R�Ipٲ�{;sV�>Q_:�qr_Bd�#�`t�˯�ˎ�Ը���&;9��� �Ǔ�l�R�~�i�[��0�޽��Ž(�HS�iIU�a��>ҎH�!������3�+5��>%w�?�u�Ah�Em��C��՚�կ@
d����q���-ug���p���S�!�O;�{}%���+W2� ���U���J`��"�����?!�3U�'�o�F�:�����q���]I��,���4z�3�o���&c�Å��i�3on����	��7���r6�ȃZ ��R��ño/.�ūR�t���DX�N.8cz�}��K�upac�:��쐖�ΩT]-���=	)iP�m{lJq���X���j���T���d{uNee����I�[�
���A"j8�7&�Ǣ�	]k����m]j�	��j�yf�pl��B�j�ʜV);o=�P���		r|Z1����H��7y2JZQ/D+�_3�]�c�|�	�Z�r�q�w�(lnp��)FU.��hɤ|�U�H=��N{g}�y�{�ΫU���g]�3�?{��?������JO�T=3����Xi��5���X�.��V�8�w�w��rx��濐�AL%)�L�e��<����i�ӤQ��������J,8|x��dV�j̈́B���ao��;N�� d���q��^Z�<~�,d�yη�=�#��������O����LK�r�a��~���@;_NPh�0���/���G`nǯ���o+.�վ�bwQl��	�A�Wm�lw�����w�N��^��,GRfx~5	��}Qq^�K�*�խ[5�p������<�a1����&=�G�ߺ���W|O�D��
�4��5��|| ���`��e�3�I�>E�|Tb��7P�z���L'�;���<>��FF��+���;U��s�4\�z�й�v�/�Uu�T^2���ۗ4��e���45��-���I�a�h����Aw��hӷL�E`�c�	3���f���#7���C��'3t�h�E���A�3��Ju��p��Fff|�!h�:�t8sQ�@6���Do��mڠ����/��x����񂩡�
o~��G����2�w��y����η�(cF�����Ԁ����u������(??Pê�(�e�znk8�~����8h���E�S,��ţO.����P�
���PqR�0��-�� ���:D�O���wN����S��у�g��1gGeĉˋ��'�E4�*��O�g�ɿ�	���7�P��o>�A��⻊8��9ˬ���-����ԙ���[,�/2x�+z�w���ʑ
���
�[�I8&蒵��Tۃ=�����9��r�{���2;:�j窴o�����S�*6�|�\-�Ho�[�A*�$�d�Q��I%
�����z����:��om�c�!�R��B�Ӵj�����tߴ�éO�z/��9��vs�a���A�j�Hc���nH�a�����Rs��U��|��Xoh~�r��I��s��0�}�2��(S� �A��yo�T7�����=t1f<�Ϗ�b��`Yƻ�h���F8���졏���g�_�-[�x�m7-��ք�7ڥE�@˴��2�` ߎ���O^�I#AI���Y�Q�@�곐�y/5���[�o\n�2Q@��k���3�e#�����U��"�g�Y�v6:+*�gI�F��7?9�(#�	*k�hWhUn	u���$���>Ji]ڋo��� J�oΓ)����:��69�Q�m=���h�7��["��{=Q�\�Z�.�*X���<=���L���Zk��B_a����}�T�}H[��.'L�L&�����2}���Ƙ�L~�ylf�E/�mkP
����M0�4MP���y	�G�^	)�F�z_�Ð�I"p�e�s��P�_�.�;MC�!\l�ǡ���������S�wn^Wv�֗WCN�PD>�x�O�#��O ����SG��7�։B�;�g���w�u=�?��Z�hK����=�򾙙��^.`-��������/D�88�f��8���7.����❶z�ځ� �}�c�Z��X���s�mD���@@�iQ;��F,�;2��͢�<�{���굜����Ǎ���ߊ���*9J�غ˷�&+=z�kΈi&��2`52�+�y��|��������0�Dk2T�]-��\��V�C$��O2�o�����@���ږ�OJ�9��|���zM��x��Z3�+��� �xH�^����}��ί�iGcj��3�d�7�Aj�R�ߵ���pf�fO�mͳ�%�R�]�X�C�d�@aO̹�UIv�,LE��"�c!�q���/�M��a�ψUj�#-}��԰^�l���@,���B����`��X���9�s# |v�m+l�|ߝO�a��ð��Y������_γ@�f�7,��<8\�c���kH���'s��yCѢSr��D��M�[�:�+`��u��/6=(�X�AbB�7�GD���Sr�M�`������״��*�/(Gt44��{���s�z���2���Y�&/�EƼV���˔��1�¦M���	��-�:.9*�!�]�
f���jij�U�s�u�s >�*���))���st{:�8S����	������&��Zܹ�T���[�
��D���qo�8S���N/��:;�cF�2^��!S��۫W3⍱4�ls�-Z��&�,����Cm�%������\���r�_3 |���.y�����y�*y��� �*/�w�������4)�!�O&o=0m���+ǆ\����:/^��P௦%CQ���TH`���D��oin��N󩡕v���W����z�;��D��tF��
�SQ���R%U��>L)t��>��HGWc�4ßz�8��I�⸳� ��O�#�q?�g[э��QM����<e�g����͉�+dAڼS�T��L֎;�4��������30`9�����#����{7(}�2������M&*W��x��BÌ,����&����O��.,�XJFE� ��;��+'�w�(��Ի��c/?����Q����\�w�/A����
f#�1أL��ظ+n<K{�7"�<���K��2.*r^񻻄쿛�)t֪��`���v2�"���U�5#��,�.q�6�-P�+�**��_?��<6�l�
��K��+E�S@�;�=܏|�J�r7��J��W���U������Y�.fJ֖�R�ܥ?��Pz��E��*���l$ �t�-@���ǨEj��(/����y{22�����Q?�mK|X��\'sQޟ�`�?�S����>z�q��D_��&z��z�_�.�G�o<��֜u4�Ǒ-�Gb��hV��9+�(;GK|p��7�� �9�C3�7���.��-��p�|��t���f�<)�4'�8�]�jqb����D���C��0��%�4n���4��O���#�9�$Y��6��N$���S�Ve{М�<2%��&��v�\�˓�Y�"3�j�S��?���L�p��	����:��{�%ΖI��e0{���x���I	%ķ�;p�|8i��f���VwBG�����QQ��4y�S\�{̦���ֺW$7J����N���4i��i�9�!3Y���&�� �E��q���yX���H����>� L.%T��Wϛ�Pd4b�oX�_z� ��Ðm�����r�*�m������\�h���� TO?�����S!�cGٛ�u�٘����4��q�lw�>�4�W.վZ�\��)(��f�vZT=�R������C��N�m��T��Mf[���K�`Z��q�]���Ch�*�,���r�j9R���4��(d�Ho]~;ѝ��2bQ�M�Tՙ�JyS���u"�?	��b�ђY&���^V��f@�Cixtc���M�0;�����ZD�sWg����j�{x��^�(.�ei���?�������Ǿl?�R�:́�'X�>˂=�)~�i�{�\�^�X�>3|�AIQɲ��/L"go�\Q!�� V��������:���,.����J�


!�9�m-sz�FV^/�憖i�ЊR�ߴ�=�2#��d�?����� ��� \p���Ħ/�8����I%�s >���ǳ�a�ue竀"��m�ɳ_���U��,+�8`���X����k���č�[�rLr'�:/[�)G���h�3�/7�%�����g�5��?�쿼?�?�����M��8;V�S�*���*`�^�4��<N`o��R1�����rAG�����&_ݏ%]����C�%�_��(���z��)ѭ<J�Wll��w��2MSnb�±1��Ɵ�o��0Kk���E�Wv���FQ�e���>z����Y�0���� Wz��8�ښ?-�8=��tF���k-'�8���!��	q��V]t<�&�u�4���-�g��^������=�ۣ�����
E�۴�����e���LP `��r3��^eIgk̀����L54��|;���������.oݓIH\-�4i�6DU�i1~`����ƍ����,��	x?��[�Q�[��6�Ƈ��]X__8�WFn��+	d'9�XX ݴ.JA��Q��Cy��i�@
�;���N����b�asDcW�U�N��z����/q��:V�X�tj�(ک􇢑�_FPm$��qu#+nT�
�ޞb�	�J��|�Ţ����a�/o��K�ϛ)�Pc㎏�=�0�gt�$HG����%1q���?�����;��V��k�b�2���K�n��DU��S)dr�ySտ�D>4�pW�ߨU6o�sY>[�*������g-�lq`�n�"mE=�=9渢�A4U�l�.�|7};�=S����`�=���L]��呐@��)�������Uo_���uR�:�P���|y�Z8UU�o��3�Vd���{�7ب���6��,��-S���(�i�ҋb�nqUNٛV�u�:�kpK�4l2���{�[A���Ӭ���k�Q��KE�Q̑���:N�VRWqs�:��U��h6_�Q�	x�G�0�V��롡�/b$#(a�mn�� kI�gR�bmC+E�u�*��i�2��t#R�	�[),��\b�l��B��?���I��9/���h�K�!!V�ʱ���W�ATG��B�?p%i�
�F-�(�*�H҅Je&8�� �5���07���t0���c��&�EY��<g��N����"�_�<ٝF�VV�hՖ��������?�k�ywl|� �<��1ʸ8V�	ĕ��i�+zi��&%�QO������#w��G��@�ΎJF tF�L�TrpP��B�C�z�7��[���ŵ��-�~�lR��Ɍ����<Xf���BAAy��65�H��{GtC�+=C��Mǽk*Q��L�땅�[q,u� gh��d!5�Q����$��w/��I5=u���i����$���H�[H��r�q�
��F3�}�h䯳َдQNr��.��e��Ph�l1���8��q'��
�uD����l̆�M����	�ˮn>��ET��D�A��)#~ڵ�y��z&�>ݢ˛2b%�L��6�q'�����癝y�O��_ˮ��wH�5G?�Jܽj�v�B�5J&W��2��a�R��0��,q�XF��y�
��`e�X��G�O��Ú����y�ӧ�x�<"�b_E�X��#.̆��Z,g_]�PH�����U�~.�;��/��,:��S#'R�&�WH�%��؋e�Y,�1�$�aŹ\�Je( �p���3��������X��w���}=u7�ׂ�ǃL��rO��mMG߇[j�2JeĊ
3NBo��
���~Qnv�<��W���ˏMA{��Hu,)���n:h,ޘȟA<$��8=ߨ�+ܬՓ��ֻ:9��0$�R=��@��X_��ʏ�<G��������Օ���g��t�����hE�㮖p	��y��Q����Ɔ��	ݹ�:�����tA�Ck}���['��u��;�%�e��N�����4@8�8G�Ռ�ޅ@ ����˯fXc�6���@7�ӳD������H{;o�I�h��<�hg/1k�Z����ΰ83�V�O�F��áK|�	ࣧ��L0kX�r�H�����t�nfZE��(;g���lvq��X��v���x��v�'�?TQx��HGE�2���h�[g��Rb]sz"�����@XT���-�y���Xl:\�;�4�l���'�#�j�v�\Q|���b_"��a����"�9]#�?F���NR�וm�����io��7u�u�`��_�0������� n�"��W���u��T?�H,��گ�惣RҎF9e�~�L�P�-���rXi�j�R=�� ^�V�����pH&���N�'P׀����=�)(��w����vC�S���el>>�ph�;�+y
�q��V0�]GsXⱨY���m����Y���U�U���������t�Bͳ�� }�+�O?g���d}Oz������@�L
2��E�E���g_�]�,�O���f��+�8���
u��+�邪˛��#�ʢX�I�lΰ��d�F��{��Ԟ7P��.�D���9I[� L
��m�`�X��#�7H�K�8�$��2
䮣�����,k�g�ⷣ��T������$A��p�\�Z������Ŧ��bv���`�sy�&�y\���^X�Q?[Br��/�	��g��&��}���&[(HεAN�iTq�-S��aw�.+��^a9D�_~��L�p�����:J�<jq��A> n�f"n��X0�,	��5Cl�1�P1N1��]H+���?�U)�K��1������9�s��X5SLė�|Q��g����Y�3����%0�%�~�z�E7;~��<D8���?-U%�V9��s�����_3@K&�����u�%�Rʆ�UP��<��Fq��;�oUڏ�N�����ٮ�tm��������C��ʽ:�}&�T%m�; o�Э��KT��JqD�ܾ@�b�[t
#I�)?�sq)AF��)�D|o��S���]`P��+LK�,�1]�FF2@�I�q��fv4<��41]Yc��F=(�@ξ�,"��t�ڬvM�5�وᝥ�T�S�3f�;�W���;7_~6�[aBo��%�?Q���L/N21��f>��.w��#��-R�E���?K�o���� �������o�/�Z�z9s��}2R)���{��9{`� �]H{U�p&��zN��,V����o��(I�#���_9	2�v@�rv�2����^���	�:��b��i��Α��0~�?����]���D	�����A�Ԃͅ��[�$�t�X]}��7��%l��P��pXЪ��w��Fo��8pIE��:0�$:��n�̣�d�OL� La�y6u�`��Q���ƬRbbd��8��[��DoM�Ċ�E5=D;������.:��ʘy��΍�Y�=s]R�zk��dT��.P"dן��h�+aX�
PMv��r�&��TzmP�5'^qc1�����	5&e��j��W�ƛG���;��c(\�CPm�t�i�Qӡ�W�kM;;�R5N�7<v=k#�@��t)M{�R"S�\/�����J���f�z��܈4�-_jh8:{���љ�f�x�/�D.���ܳ�� ^�i�z����~�B���'h&�kq��7r�������Qm�*]\�u�Kvp��Z�����cS�ݮ�5�v}�o�c����rY���@�������J������R�d��Z�$����H��6~uqi���"���t9�B:I�3f/���� }�W��q��H�,��FՓ�n͖�&}W�[X$�*�+/�N�.���M�Ǚٸz��<�~���b]|6U]K��m�� � k�QIK�u���29h�M�LK;Z�/Q�Zh��|�:�ȳ6MG2u�h��o�>#��<g56f�:�rݨ�c;�~��͜q��a�����z/��]��6��6�L>bӌ��FB� ���Fw�wv����ã�������/�2}�yF7�5W>PR^���r��I�
qtO�zv��4�ڨ��0�X��p9pko�X����.$'�L���x���g���*Hݏ%Б��|�I�>9�;���K��bو�@hBm���V�?ۗ{0����ҫ�84�LUpӋD�+�2ρ�w����~$��1��k^p.=�˼���ϙ�����+o�FS����۬��z9Ѱ놖^bRm����p2�ʁ�����#�с嫫��'n�z�a0��]4����p0��w3mu��4!�ƪ+���	���	���~#���Z~�WV���� �U��҄m�IRq�W��� �=>�:�e"�=�Y-b1�w%��; ���A��ہ���6P�6��(�M?Í�m-n�h�Z4���O���,���n!�釤��l�o>#OЛ��`���%��Rx���CK^.�6]F5V��0�\	-�d�On ��	=�,F/g���a/DlZ����Ӷu��M���E����|H�M�zB��#���+��Fo�ԯ�gMr�nN��-G%�cv�1`)��&���.���;!r+��ɽ޵_;v��1����p������z:����bo?��f�,�`�^�T�ׁ�W4Ue�
�4�=��
�u�#�cs���((<�Å�v�a���t���8ǈ*SI� �F��8�ԇ�����FS�����m�vFVo������UW:|�����{&ǵ��ݰ��6�-�yZ�=Ű���#+�߰d�F;r[�)��v=��M�H'�=	��
{�ظ��g S\\� ��P�A�-2]4���B�MU�1�;1n*�!����f&J��^�N��1�E��֮��!�����"�� {����qz�S��!�oY)�>�{H���o&��&�S!%����2إp>'!km]��?"�_���g���:��sG��'2ω��W
����Y���C8�E�l��>��)�i���O���,\#Y3*Q��U4�c��kE}^~����מ���(�)�1�vLק���n.��==Y��Ԋ���675��d��(b��|�?�a'0� �(,3��2�'���I<F�%�d׶f�-d#m=~��`F��q�xIh�D�����)🪼�J�̉����;Tuy��y�\3g�"R�2In��%5aI�+f½ޢl�t��Y���ڽ#ʛ2��Ŋ��2��A<*��I8��eD��$��J�q�Z��pjM!�LA3�K�-���y���0�V��F�$T ���h�H�HW^��N�\kĹG��^Gz��:�~�ac�����LM�CI*��zߐX!Ϛ`F �N�[�N�+�^�	��;�x��a�������q�w�c�Ʃd ��ew�,/��[��䷌.�ar:B�u�� �># �mA����&�������.��៯}>����CQZ��O�^��[[}��0���g�kY���ǆ׼���*��*�|�ɰ;8�j��׬�?��Ĩ;�����H�xsjD��ɵn�`�-dў���kg�2�{l�U����L��{���:��b8�hsB_9_���'�M-��MM�9^6 �.j�H�D�D���61\HM�����vv4�uM�%\6�}��V���Í�<?�rS�Nғ���px~��H��~�u�L���u���� ���U�h�{�%��yl�!{߻��YNGҐ�4�w��M<����d��*��lle�d�`��D�7�Ɲ㢜f��WB���J�����O,z)�}9躌�`�k��o���>U�g{6�@H���1��o����#�<��Ŏ�Ђ�!��^*-�-��������hL�8��w\�޴��t�cJ���{~|�W�	���x�+}��C]��8�w����uz�Q��D�̇����������J�љ
�qP?H��2N���9	��o��ut6�)(�h�2��Q�\���v5�徆�y)9�th|����ȷ�B�D�j��ğ؊!M�R�U�^S�7`�����Z|��N��<�����p���u�3-S�0X�Ne���gj,���r����0c��MU���/�j-�EP\����E�X�WKS	������ ����LrXCDq��[�8k��/D2��$����m�< �Wz����Zn��JI��d��棶����6�o��;��U|@$�����t^{_`ڧ�}��Ua�)��� NU�1�j�Y�7��P:�/�S%�t]5q�6���E�Z��b�&R����DCRuUOT�i0AL�C�x=I��.X�s;�����Xt�ǂBQ�c�T/3�.j�'oWk�o V��W���:{�n�~ƈ����e���-_`ܭ��p��Ci��b�n��ݷ��w��o�#�3�A7�N��,ŕ���3�uc�s���T� ���q=��2�7��/�1m�kOؼhhQ�0��F��Q-����O4H��s���~Y��~�Y^Z��&y~aw�6�)˾y�6��m��`����_�����m���y�e��70F��y�˙�UXR�_���ym@/�c;�&⣪>�LM��x#�������Z89���.�
 c./��O���iڟ���έ�� ����1����� j��$Z��-|�*�-63���L�g���:�P�G�a��n�w>��-x��i#���Y���Px;�)���nIy���y��7h��C�\�L���3�a0Q=�-$�d`��,D�WX�W7��ì���{���?)/�(H8��>"b�K����'�ט;�W�G�"SL�E�R	 ۼ 0
Ў�>I�ڔM������ӥ�;��i�սt�Sjtr�6x:���a���D�k9��?�{���7�o|�XgE�?�B��3�BL���������m��;���WQu�N[?���o-K,}/�1G��AK�6r��ʮ�ۃt�K4*l� �]i�w�����8�w~m�:�� ��ra�j���_Y��[����v���eΊ�¤��I�NTq(Y�����Ǥ�	ٙ\�/>t���&u��*�c��;�@���Թ���D��]!v�3�4�LO�~��p��Wh���lB��e~]";};a`<8�޳B@���(S�1�0Xߗ���;C�๽/\��L���ؑ�bb�2$y��Z�"�-�t�[�-���i[V�c�bV�Ox��1�{�׀Q�&��g�rbSD<�R�;_�j�bt��|�5a	��o[D����'�Gg�F�o}os��K�W�~rd) 8!���z?/:cV�����;?�ؘ"{��`nU�0�I"?��=,�!i��]��L����Ӄ2���J�=5! w�A�%�HQ�/�����km�,^����jZ�P�nt�S���n!63ÿ���?LO���	\l�O@�R�����)h�&AM�5��.��*O��~���k��B�XV���1�y������Ʊl�������*�G���������;�y9�f ��|��E_s�������O��˒���8�w@�3�ƻq=�\��&������,�uyiR8��A�8|m�v��I��wC�_��mI�,60�]��W�0��� S�3�`z�թ�h/�P5�ԥ��'��;;��a�>����4�����5:�8�m�O4�����v�Lg�y: �	J���?<�`3��Ȝ�8ɹ!U�zսa���܀���X�1����D���|#�G�YT�{E߮�f�o�f(� -�����NDX�c���Bp�Xܯ�qK��OM�0S>��1qI�@ �:��REB� ���s�)�r��/���*
�'��#ɹ��=?�E�&�{I���9�y�P+*�*z>�X������a�{���?�5�1�	fC��4�wR��ԉ%��į�FW64|�мK������!��p��gj3/�b�,�r��'?���'xZ��`W�
:=�у�y^�����1T���nQ��i�1b��rx��Pf����?Q�Ȝ��fs�OwN���VG�[��'1���T�!����6얿�n����Y�uGYY�3t��0���ݪ���r2�ӭ�,�Ǜ�.�#��Ӵ���8����� i:�茞�iJ�3O�z�č�e�Ԛ����OVw��fL�tT�k����=y���jd�;	v�UI�s?dZH��T?�.��x��b]��`�i���y6�g���;���׳ W�Z�h��SW�$Ժ���>5�K��1axw�20�R8�C�T�Ծ�v�5�e`�pa2�.���X�J;!0!�h=�Hm�Zr=�,5LQ��LEv[����xm}1ѵ���a���Z��2���ؒ�{�0�� um�«�4���'�}dk鞐؞xv<i��sJ�ݬa��J��F^��-[�<ŋPQ
��8�~�]�@E%�S���NL�t��ܧg�.��/e�?U��~�qH_Q��O�F�S�#N`4mA'���}I��F�=G���B^�Q򗺔�L�cQ�<�U*��(ں�qK�q���^���m����6c���� �ȍ"�{��)}������XR\S�yɄm8��`�o��<�؋S���I>���X�i�}�b���Bz�e�&�,[]�~Ɠ\���T2`=�(�O�I=W�(�~8.�V�"n��R����4z���~��T9�Z�In����f�E�/���h1�2z	ZC&2��=���L�����t������U����w�,t&���tz����{��mlU�T�l��>�c;ޛ�Q�u�;<�.�=NNM�sV�����-�׈�<�+�t�C�h���2�I�h��U�G��	��~OL�B��3�IJ�h����{�yQڤ�&��l�J������ܨئ��dhi�OW���z�y�uE˟Y��moo_|cJ`�~�s=�*�S�#�M�����q�@^6�څ�~���xi���.�k6s��gG�3>z�*��+�8�v;�|���g5��N��ݭ~��(6ARo����3��A���l���"x���AJ������-�2����"ûw] ��Ú��y�'��4�A��o(d}\��!���93�<҂ꨱV����M�%A;J��1�����������fW��v� >#��x��#,s`ذ�N�X^�Y�:���4%>Û��;�JuY��r�h�����L�%	4b�/�fL��t�*#�n2�?�&���p����+�q��sX�F��;%$Xw�]g�;Ꞝy���ļ���C�nq'i(�����3�R��r8X4h�r=�Wɍ��8�
}C�q*�CE��Fc4�p���,r��v	H ^�g|�az�O�k��M���,��`�Fj����S��>?%�� $4�A
�x�Ĝѻ�������@ Ս=ÄÝ��]��� ��ύ�5QH1���1�cń�GQ@@>Z�A��N:��>PJ�80�n�P4JZ��R\>�s�>�j4����=��ϯD�h��!O��btC�w�����΋������vz앤+��/�������n�{���<m���s����3�Y��?���˳p�e�����Q�r{����r��u���6׏B&�zy`z��;+&��ɶ'�s���� `�l-���)*@�8(�Mo�Y)Π�Q�Гǿ��0L��Ks�D�� �	
�Os��^��1����1�1�� jvG2��������3)�h�A��V�F+司�gd��ߟ���aN%3���h�߫��!o!��
�������K\1���s�A_�%N�8���^��S�/$m8�u<�Ӏo?��lOR2�Q����	��B�m紐z�j[�W�D�<3[g�o�N\z����:»}z�J��(V��s0�L..͛Ԕ���{���w���幨��Tw�����VSII���H�im���m� H�Ԣ������sN��ȕ�[�Ȭ�E�d��_�!\��4 �����Q�F�W�&R�ё�9:��p"GC6�8{��uT3{���s�_73;�����<ڲ*�#6��&#&%��,��9k��Gh��J��[;*+/ϺU7�r�<�!5�z���*w��ɏ�JX��dqY�Uֵ���.�P�b����(�dX�i_���*鋪[y1;g�_�_���>S�Rë�������:�b�w�ѵz�=Ձ��;�I�-�����s�&�?�Kj�{'���P]V��tb��X	Awص�*l���:�X��_�9)�����x'����츒�;z��� �������+����Ԛ�|E-hm�uyVBw��>��7XYO������=�}t�c�J_�7���5�	��� Sڟyb�4^G$�<���:,�'���g��o�< �]:�Jh7�����d��cD���Fި&���aŦ8cF�5e�B����Y���ڪ��;�Ν���w��C/�o�����N ����a��*)����4���)������t`� �@�R�H�"?�߳Ga�Q��V����V�����?B��&�6t-Uð�S-�a���b��=f��]��V�-m�T���~x8#��u��¥�^���KA>�����nͶ2yz�⠚�,O���:� (e�g���N��q邶>)� s���/PF��adrF�h��t���za&90_��=2e�N�4V�7��h�l�SS��%�?���U��-�*��<��}ձ`���d��ʀ���Kvm��$	��~0@� o���]�(�d3�R%ެђޜ����_kcdݣ���w�[��)j���29�r"������X�=" 
�'�
 ��ݘ���72("\Ec��H��
���˺{�����r`�8��j���r/��NB@O���۸-�{�[Y\�
����-J�4#1��=l��ž���@N�o�8��y�6'�������*H������7��������%�ކ���J	�Y`�����6
?������0&�<�q�9�=)���Cr}xe������1,:���E�����m���P�cI�0�����a�nI��驖E!S�B�����L[!�y��wj�	��P]4�'�\�?D�J� C_�������k����k�l :���v���j��\D �9ڙL���m�S�+g��W�� al�����N��M��%��{V�'�Nz:�h"R}�|�ި�:���-O�>ŀ�#Ex��OC����g�;5fO�,��Q&���.qN"<�D���
~���<�閤��D����,|+�)�sM&r�s�rNm������~����]✧���{y�����R懅@(�!��W�	�#���~�kZ
�Ӑ���l���_�G�Mp�>F�ptS\++緆4~������\� w֔��n��?j�""WF�L�Z�B�7�G�A��_�h�s���Ua���dz�^"O
w�?��_Z')��7�������]g�y�-��qY9��V4�W̎�=�p �­Z�M�A-�*��"�+������:�-}j9;�R��s� C�\h����46�o�3��B3=|�B�5lD��i�5��`��5��Մ?��߲��>ݹ����J>H�yt9O= �	�-���������J���1�Q��1��R cڲw��μ!:g��^!,j}�A����g���K4�i��eb�Y�y��'A��4������� au8�2�mE�v:J��o/u5z�{���oĻwn�{~45q^��|�,�&�_�%	uo�F�{�i��fE���`��D2�6c�,��8�K��梈W�Q�(c���"B�<aG0�SW��#w���c�Q񦑂���T��e��=��̓��M���TnjJ��c������?����4�j�"�a�ϞȞX]q�7���E��K���M]�b��m�Ҏ'�o��|��6`�mfl68����	�턮��Z��������v׻���x)���u�����Ǧ�U���je��,���f�N�%,�?�`B��ܗ�n�H-]ݦ��
^ދ�B�{�]�Phpj����\��49M��P��Q�-/�����!#B�oe�U�(��D�NT����c>2��i�N䜵e�W��O���p��H�|���GQ.'q�MA=�]�5vm<� `���l|�}������T��~���{��A���J�b�Y�v�I8/q�3��Q����x����2�gՐ�X�G��`�Lh��!M�����S��v�Wٽ�����N�j������>�/C��R]�\"('LCB�=��=��׽�B��e̐M����ۧm<�����]|��u��m����}�����?pqׂ�F��"�g=��E��v�we-{��E �g�YŴ����}���!���x���{KbM�8��oGUf�x:�7�JKX2O�<'�X�c� ^��8����Փ�w�c��F�q��&��>��Xv��[�����
5�����_�Wm�����Á|*RhSi=M��\B�)� y9eUе3�-d|����̟+Ii���hG���V��"ӫI�yO�1��I��m�t^n'�����:Ϙ8]�/A�׎F�(T�9�,v��퟉�K��>%���?�Pc= m?�G� ���z�<T<Ll������� ��c� xӥA慄��p����=�!�����,���^���˳ӱ���0 -����fڣ�uġ�U�8@sN��s�f���@�t��uP����Z����H8��=��Z���ከV���v��#����Ώ�N>��:���#��	��*���7�S4��X,��P�R������o-�"M�陸��M!Sg|���g.�|"SJ�����{̣�o<���01@!�_G���A���rG�����W�5�5�ߌ�����A��ng��nz8�߇��ޞ�����D�7B����k=�!K1Ւ�����G[�����(q���*nV�r��Lq,]^z�:��b��U�Ou��OK%��̊(B��J��^]�=.½r͆���{�˵�����ƽds�{��.��������#�z�s���x��9�Xၗ�q�d��O��hCN������$�U�pU{�~�O__T�/F,�O�1O��\�r8������������e-��[��U��K�g��+p���o����@h;D|�����y�=�QVT��`~�[q��x�U�Nk�����@��F��T��K#@0��|7��c>^�i��sV�؈7���x�s��a�����ms��F������Z�a����ue{&%�jk����jC1��}m�eu�φ�ϱ�pwƛ�;4~Gڟ|��h_;V��<l�j�.���q�:���0����s<�oӰGf.Yŕ��e$������_EfoZ����֮�TS�T�⡎�\pQe��)�H���9y���Z�z#�ț���G�̦;�I}��(V�%S�:g�&5�	F�M����-}y06�6�?�E%���H*�d��_50�%?��2z����I�T�1+S���Tѥgѫkz^P����=��*@m$
�y�UP���Q%����,=~�X�Q�J�Cmߒ�����/֊ѭ��x����N�E]��@�N��z�l}��R�9.E�K����O���$�m�
q�I���T�}J��J������@,)��R�.�[&vq ��V�ðbp|��EK�r5Vr�9��}p���G�dQ磌þlx��C�A�
P��+/��G2_�dXX�'����w� %��S�F�S��#�3O�~��za[;A�؛��.�6��P��َ�{��y�Of 8�&���EO�_��L͈fM�/�N��l�UA��8���b��mI�Cᄾ����r���q���S��.4�&�l76�;�4y4�E
%' g�C�� �����nBR}%A���ˎC�T��-�7<Tq�|�L"��?Τ�.?RXW��*:QQ(q��O��&��-{Ќ�&W�h��̃�F$��}�K��W��l!�P����$�2�ܡ��#�ϰ�������G��Qf� ZI�~
IK�=�(_������
v�6%�a��(?�:�I�-&,5u���l�K�tI�U`���Owp�|�NK�i�M���a&,���l}��^�<Nɭӽ,+�ƹ'/,FK�M>��\z7Əc�p�taܸ�VP&�B�OWZ{'{a|#�D�չqC~�<��޷s���� �.{9���T�Y���J�!r5'm�����ȥ9.��XhN�1	x���g}W���/>ICii���'8ܵ�<B��i������v�:��xp ��x���1������a�m:f�v)BEB���{|��O�	c�~lJL�?G��9��^��<�R`���k_aL'ka��t)1�Ȅ�%���8���`D�ŠԷ��\�I�9R�	ժ�񬙮�\�jU�*w�$ٰ�QUޜ�ո�F��}�$g3��>8ף}��V�4K�Kes��'=^�*�T[p�����Q�I�Ӥ�e!�S=J�`���50�=L�`��$j��7V�)He�1�KM>F�>2+�9<���.�c�v�� ʁZq|\��[[�n.�����%QQs��\�N�M��QKK"��"�r�'��������NL��Y��^���x�;���I���a��*���Iyff���uM!Tg�ew�G։�§#���M"������ �QW��)~�\N��q�Z��9խ�?9n
����ɾx1��S{G_S @+]�X����`��Y�h!q
���C���^�D�.}_�p�#G2�]aTU�h�i�l�������'��["c���3f[s�=_���4����N�����[h��T,��f �4��s=��r.�fIZ�:��~\������C����~I9�^��N�^��xP��q�ظ]��Ա�L(8q[S��y��Pw�i�)������r�w#dS\����oB�>4�'7E�$gO�o�y�dZ�}�s��m�\m2)��7�;Mɻ������7_8騠��>	�C�І#��wh?�Qv>mu���^\�#�*�������Ċ_P.yqݳ� &곟A/+����ؕ`�uX�������d�B�~�1�dV��c�}rV�.}{��.`|x��(+Ro{�
�\~��^9ldW�Ə�"��|��n��M������*U�|,���ۊ$N��9��*,{������`��4�V!�c՗��4���_�5��Yu��\�1k�\�7�i"@�[]�n3&_W��5�i��2��`͚���\�^��
\�]){2n~Y����MW\���NNsH��S��f�\yŵ_���n�&�L����;y�,���2/.��u�{�k��c��`��`]B{p��VB}��=�esCo[. ��ql��'�!� $��l,&�Rř#sv���n��Y��#<�;F��]k��� *�z�i)�I��o�Y��`����#�̎N�|���t����E=8@����q��H(��Я���KǊGtƓ��<\�Sp�x�Kúi�$��=
%��4�(�� ��6VD�I��o�*�6L���Z��nmѭ�d6ޞF�!u��R��G�r:�Y�'{�B>�`"�W�Rḩ�>"�P�����p��h�����&,GTq��}F�s�< �<b�,o���14=k�o_r�<UI��!%©^�� �?�R�=�g˼�rp5ZӲ�]��Γ�!�U0cc}9��S�v���i�M�rTԲ#������;ibu�AS���Dx�����[J��d!�g�����e.��N}8v@ ���>�o�"�=� g:��{�&>��E���iݏj�^��^�t���)�jh�P􄉞�kx�O�1�8��Q�ޞIm][P��ƍV�	j+��I]>�eOYQ+�zajs]�x[$8sn�C� �؃{و�p������Z���cn�L&�(�5������~�cQ���kG�[b�g��}�T�{��/�.��ͥ���m�*ƺ�_}]C�k�.��G\�Y���kF7K���z�]j0v�T��Xr�̭�]����1G���-BF��b��Ԏ֎�~�Vr:���c���f� c"��Y����߮
��Y��������іvKn��:��[���䫚�h����wFY�}�ǟ�ӲF_�����4L�!�^&�����_����+�'��fWސ�]�ַ��4�B�A�����ʵ����|�k�ۧ�{z��=%���*2`*eS�|3c�>E�j1/���'l��X�^��1�o�o,z	���'V�m�֕N�/��� �����A���}YZ-輳��-tl���_�l�^�t�8�l|�d��c� 3	J�����U�������Fd-���ɗixDZ� ��m��RA#�R&v����a��~X�����.�D/���n~V32��?eU���(��2Q޴���]�>�9��j��>P_1��� �Aյ�I�[��ph�su�Z��1���Ҭ������"5�0p�d?u�<]
jɔ�:!i��GNqZ\z�:�6���������Kn�F�����J���p�����F$F��:j�8��em��0�b���+"�O+��IB����s;A���ݽ���9f~V�곊�2��F����A�D n5����y����7Uc<K����y{KY+9��Y<.��"�A����X)�9y�k ��:j���)�������:W�x�nU����Dl�h������NЈ��>=HӲ����N��y�s�����"�.��������km]D��#���9/TO�ƺ���F*�S78ؘ�^��2w���'�N�?	�υ�FR3C���)��O�z;�T�ׅ��,=�
�P�攜�;W�K�m�)������������ތK�i��$!���Ŭ�D��~�;6�q�,��뜺�U+�q�/S�]���E�x�8��/;~y$r��E��?I��}{�cX���Vea^0�	Rz�cS!�&�>��C�\����ڗ��u����~1�JSH�5�ܔu���0����v�XP��	r�-������/���uHNQ�yhaۍ�+V�bι��U�m7��NF��� ܝ��x��5B�o�s�Ӣܷ�! �G]�m�^\��'&�@Ta��p�?mE�8jQ��dH~�ɷc�4 �õZ�,B��4���5�Q)o�Ld1Y�l���������oKdk�.cJҚv����^Y+u�ԫa�l�X5��H(��
kƄBI�_�/��Y�����bAV����Co��/���6�0� B��2�:�n�䦮�>bjm/��op��P��v��1�(L�:�ݘۉ��Ұf�Q�d4Ã�k:q��ɞ%����Yx�]�j��]�`���tr!?w�E��Ԥ&zkmDʘ��p;>&�H'�^YFBi�{�&V�|K���(|��Q��߰O��e���PQ�C�6oԦ��]����|S�j���a������V�F��b�O�&���qE�r�B��"{�T�C޹�Q���Ԏ]�Ժ��e�R�����W�0���������ϔ�"I�<u��:ĺ�%���#>^��c�V����X���Y�2��ad��*���/��-������ �s`^��NB=q�o7�79ʽdH���"��v'�i���l�KI�e��2����MZ���?�P�]ߖk:9ř�X;��!o�p��X���nA�U���C�mR
7���I�~3��HU�E�����A_i��W&,��l�ߠ�o���lt�B��ia\�L���}&h��a�� �	���Oh��$D6�3�2ƴ�4��7�;�3�,��tu[��G+9����eZ�o�����>}��Ԓ�$�Տ��#����'�d���oK@o-������zi�����i+n���`K�Q�I�WGՃC�>�O�ڍL���Յ��	����8-�[obC�$��)�'�r���1ﯞ��2�Z�FՂ���uN+��y�x�Bi�nH&P�y�T,���m^Ndg���c�uXI�Ze 0�ҽ�5�Qsz��ɐ�8/o<!�h�*�I$z}#����"��[��С�b�F�5���b�M���\���K�O*�ª���d�r�n|�I�n�^���8ZZ�@7u��z�>��}�FR�,l����%�����Kd/P�fe��>��r�=i2@�Ε<���E�?b�m��#FLs2���؃Ͳ'uo��\#s�������O�Z�0��WY�Ǒ��k�f����4�u6�����gŰ��ˆ�tP�O�P�U13�D3���/Oz�-�Ӻ��.��[��B�L5b�.�7'X|!�V�����j/}fU��9�;��# �3�\�c���3.��+�����q�M���m��:x��e�xn�;��r�hN��o΢��4"�ն�`wґJ�o~�Mp[�C��U�8@w�Y��a+��w�����s0����%�e�8Z1,���V��w?#��G*�Q|}�������9BJ`�I[]���a�c 3��u)���*�`�h
�e�W���Q��iսu�权�z%��]ڋ�a6N ��˿��2g+��,]����Ue�wN�A7���疚�b�o�}X%�:��VeA���м��m	$�E�����!�nݐ�˔t��=���Z��F�艊�2ZT�-�(����wK���?ͧ>%�F�	�DHl�VSŌ�J^��Y:���;Bk}�-������ȥgY4�c����O
%�B�N�H���Ƹ|��#����e���t�%�wΆ1rUJκn;��}1�i��
�S�� F�EL1��"�qV���aA�I��!R3+���V�����	�^��x��=��&9�҈�8숺����<���C�v�)�e�'!2�m�R�'yt�˴����\Ѱ�0��\�U����\���A�����#@�V���68�M�l}�t����9k�Sp��*�u![RRjl	;y<a��g:�2䍤��fS��g���7I��}��FOՈl�$�r`���[lL/�}YzV=
�����[6���}>t�R��ޮm�^�)�-���s�}��H}_��gQ���H��T� Gr�b1���Y�	���u��9~7/�.)7��4}xH�-2�w�3�r�Z�[��d��9�zN���� :%���1`H���&;u.�MM�� ��6���3'_�<�Wl����H���ԧ}�J���\�`Yנ"%8��9񘼊f�c#�ӟ]�`n@��or����)j�l�J�e��>b[5��W�g03,.��q�eJ��D�ݢ��F���8�<h������������=������x��e�9���qEvr�г$B�����]�="���m{��G5Я�_0z�ܗ)�P'�%�g�Ǐ#�m)�c1ߠ�)����Df/�v'g��=��+���
O������4��6�9��]��^�������h7V��L�k����.Pu-�OGKZ-ސ�H~&�Nk����g�{��4�3�ubAGA'�K�++?������d}���g�4��|^*$柭W��@�Q�����񒼰\+�X���;S ��Æ�0#�C�����e�L|��[<����g�N"�"nQ<��_�3uhV�G7̲��cbl�s�_щ�7mV�Jd�5���]JtŠP��77���ƥ�E�f)��{�^�KF�iG 0`$G�9e�m:L��������a������޺���e�X�|�,zXc:�yԓ�a����#;�)�Y^��ۚd�q��*�����h�����kT������9Q�����M>��R[-�R��z�j��#$�Kg��9Bo�֬��lV��j���٧6����yiZ�7����o�㲊��y' g�펁��e=~��ٹ�QY�����r��r��!��oW�#$%ꠄ'��ѻ���+s���H��yA���_L!�����(��,Q�҃ �g.�>1���\���4�Gjǿ�]�&訆Y��,'�@5���+��{L������eX�SM���|�#C�����޼��^���qY�;S롐��R�ց�q[������

H~��.aR��c"Rc������t�Em����a�����li�����F�+ڱ���ϧ{��E�����Ẩ+I�}z.��Pl_���1(�V��k���5"C���1͔���=��?�?��V�uY޼ruy��c}B�`D�+i�^|o*��r��_��g*��K�lu����o���ij�4���ډ����񥓁Ub�kχf�M�Qc�7n�kͺ����T�j%FztH���]e�0L�j�
�|nV�G�n���g���YN)�Z��v/T��qFkz4^�_����s�/��w����XOPBo�Q�瞿�)�qtu����\+����D�R3�����];��f�7�$�u��O5�dfT�"��|�hp~71n�����CC"A}c���ƾ��(J�G	��ج��{wtZ �A�
�����NnB�Xe��b{��O���O����I�W�,r�i�AV�g��^9��������&�k
.蕧L�p���1��{}�K�E���~��P�P!k�_�g�lQ3�Å��=����(P�U����\��~�dt�3�CBd�ab���PɃ�ǯCW�C[� �k̞���Ip,\�U=kg���3��kТ�Kr{�!��1��|E�����v{���u����E���ϗ�GO���xgS	�H(na��#�d�?Ar�i:r�@���]�;��������pL����d���Wkq.-r��]�#�Ⱦ�����}�����1�FmZ_~3�|T�9���?(�"�Lr��v꓋��9�)�l&b�;����G��mo��0�Eu��G����_{M����i~zSm�x	8�������g��XSo��ٺ����uE��(�O�6�^5����v�$��!��FX<�]�x���+ χ��Z�n����1�5x9�E����,�z� F�Ÿ�e� _r����6��\�ƿm۵�:��528C�np��b�v�g��I�*����)�pKFv��t���
�7Э�����b���S�~��J�n�/���U��/�P�|e�� ?:�6d�Oɘ�o.��uvμ�W�4�"�$m}L�+��&�^q����Nܥ�2��'×�͠�q�$���2'A�r�l�^{���'�/���C����E؃�%�6�d~	���z���jZ��ߴ��,?��{~Y��{V�J}�Oq��э_ܴǹ�5x�ӳ����X!r��{���i�]���>����q[�6���'#Y�$0ť�-�^�Yyq=l�t�r0��K�Hu������׫���V2�ӝx�лc'��7cD�M%Y���1�aEu+:��+^e�WPv�X�[����UT.M<���::-Weg�����=�O�l��w�\�O��cf�W�	p'�7O�f���G��`t��?|3,��N����I��l�������ֽ"%ZO����O���X:r���"sB�=aVA��|Y�	;���'i�K��6[��rH]�������U�V�j�}�
���EV�j5MW��.#�琀��G�F�؅n6�?��aE�`�s`�P�^��Go��33%�R�fȷ�gH�������~7�K�m��)��}~=7
��M�ֈ��][�j��n֌��ņ2��Q���`���g�*$�|�)>��/�Y� �̷�����}��Amg�7�\�}�k�a=8]ۤ�XR�{l?c����˪9;[�����3��+�i�$�V�;�_!\Fi 	���^A���ޫ��G���}�{?�@�O��7�k][]|��;�3�j�V���p�T<�u[ٯ�"�nM�@�_�r��!��cN����`����`H��w��Z��k�^�L����:.������r񷺜�གྷ������ ����Z j�j��(�jJ�w�CQ?V���л`�fJ j��A���W����]1�E1��%"����x#<��iɽo��7����_�SS��Z��U+	�4�jh���k����{���<e/���|�HJ�O�)�cObe]����qJ�:�:���j7� �NS�>c�V���׻��i���z%RlM�FY���Q�20hG���܁�S&���I���No�C��[��e�%N�*�'�	����MM����4>�� T$P���ʶs���5<J�d��w��J
�-Z[B2_¾����Z�Rﻂ�m���}�,���?�1��(�K
�o�;\,"�|Fe�$�'z��Á�t5`���qo���:�`��QK�DW+��g2��?��0���(�� h�뗜*!C����愅%���Q6�$�P�a�#��&I. �C�.��̥J�ɣ���G����E��_�/a��KS-�G8�s���ɺ};to5���r�+�n�^�:2�s�W�6��l�L�wY���+�e�:���-e*����/T8�Yb� ڇ��Ǫ������g.`j�,�s8�Z�ĵc�74ir�'9M�F��v6�h
�*\Z��~-��c��W�jD�x��+���W��^�������m�^B�RYt{e��(Hhb�Vi�B_����$�X����Q��| �����W8Σ�P�p�����tjg��N0zV���&S�B��aY,|�J��v���#�$7p`>V��_P��fS���k�8o��>�0[��a�bR��N<��W}�)J�*[�Y��%��� �{c�m��)�7m�@+��7���,|��4r=Na���h�̼�*vwbC�Umc�	����ӏ�iE?���p�V��D��YD��P�a�+���n���i����[�q�uuX>��'- MR�>���u��>���N����j����fkM=_
�y� ~b���݋��Oܽ{�m�	%�.�Y��u=2��?�J�h�?	���ŦH{]�R�|^�!0�6zĨfp��α���u�5�&;�8Kof�����8�\W�`j?sN�3�X��?�?`"���W$�S1>�#2�׵�����9 л�"�F�U�/�Y�[[�P;��H��>n�j~js�P�p����N|�V��0�Ȇ����N���h&#�(Oِ2�`7\�g����x�Dp'z/D��#�����d���`K�m�N�%/�����pFg=PT	�	;�զ�٨X���Nn���M��kr���|86�o.���;�5T@N?�~��#5'x���/�����O�?�S�iX��&᳸�B��76�O�Ғ%ɟl��Q��s_
���,P�"�Z�dh�X��o�׾gk�>��� ��{��K4��孰�Ş�1d���\O^�P,.�Ɉ_�������O�K^�
��4O�83i�h�z��O7��⦦2M6ݚ	���hz�s/�r�m�#w>t<5��M�)��T_+&�ݏ��}�*ak�{Y�.�@�t�����g�^� a���2�1�şK��'�����U�0���ᢸj
�i����˦C�r�i�����|��cfw�ߝgm����3�o�<���l��3�_-Wf�jM�b$-dx=�W�4;r=Q��4��&�t��ş6�
E�?'W}�����s��v�}=p+%����ƍ�����@&�h��?�TA- �+[$��4��!�A�	�+���Ł�jմT>�x(����+���^ݠ�U�:���M��_�4�*��$�_֗��<��t�\����Ί�2ݹ�������߿����f��J�?{�R���_���,�0M~��)�?�x�߸Ѫ�>Y5�܄b�CI�L��SEI�:\�E.��}��5f��?��ix!}0}ڪ��Υk���d�j-�>t�i��ػ;w��|o~�s��/��w���N~su�s�Ud-tn��Oc`9������8x&_)��E��T ��@Ξ�9���֊���NW��PV���!xy���Iշg�ۡ�o�<> g�P�E�2:����޶��H���?GY?tl݅�v��!ο��#�@�����S8ߖ8���Ǒ'Ʋ����<��D������#dh��B8d��Kz�n�o"ŎA�n}v��A�w�l�	e��ҟ��פ"�n�3����Z9�n�9fN켄^���/(�.�8���Q��Wt��]��4����c"nQr+������*(J����WL�+Y�Hsث��I�ӽp6�FD؅��B4��)�mf|��H�w-S��H����׌��t%��z�"�\ ��Y|���>�ѐ��;d���"y4�H�j���.z"ބ�;^�ZE��ɵ��>�?��L���:sOo5m������ݵu��3=��C�������
i��˵�MV��$FL�{�uߗ	D��#�{��ga�L�.��RJ�e���.3�{C���8oH�Ϯ��lzY�:��O�8Q]q<�+1�������g���]Ɨ9��b�7��,k�=F:l��?��u��ﶏ& �^����?bt)��"�C�|���9����wP�֜���I`C��=Y��6&*U��ȮZ�E�/,"��R�\[Z�^�QO_[+�����i��C�晃P��_H!z���)�����y����t��*M�0{$A�����p^29-�G�sz��e�4��k�!��͍��R�]P�0
鈊��������.�����k+UI�NF��찗�L�S��t%��O<�O��t�i�Wچ�� ǋ��,���%e5���p!_]��/��ܽ~�	�ʜ��2��c�wx�����of�'Z|����o�	����:ꊫ��j Lf��eeC��8�6k~w��a{
�@�О�6��^`�L(9hgH�D�/J�x�~��Ү������Xh���=��ӑ�'WAO'���ʓ����8y#O�D���{6]��~8J�j�R�>K������
p���F����-�ʃ��ì��4�U�������"��g�?Ɯ�m�r�U�� u��|�[/X����d����Rppz��P�o5�S��!��ǻXT��<�Qّ�ֹ�&Z�g�}p�:8���AY�V�TK�&)K�Խv
�ss.3��ɔJ܊���(�"&�M�-J�W���Ix~J�?��~�M���li�	�s.0˯�a�ۤ�-��{MK��|�~Y�5���K8����;�Õ�qY���G]h&���>�0e���lK��%��.��i���{."m�K��ګ�y�@/�boO���� ��?;��o��>�t�����H�$ӥ�Adì���L����/���.ڐ|c#�B��"��������~��3$�+��M�B���N?}���^�F.�4���H��K�� 'LM��������0X�8z�/M�&�!v��Z�g���%�˚{�w�ؓ�b��3p�#	q;_�D�伵͗��~;
�n-w�����ْ����u��૶�1�_z�R���H,q�;N���
4>�Ar�P?of)yt�=L�P����nt��/Ŀ�_����l�įρe�Wް����̖�V5�\Ҟ4YxK���3����uo5Uj���"���{=�8l��9�u��h���u�K�╡ȼ��b�RerP�iWf�)v2�U�<U�u�@M+��n|IK��	YH����S*���5��%�����\Z<����(&l�=+�\.b��A����;_h�%j@���E/(m�2����Y.�5S̗Eʺ��L�����8d������6�Ҳ������R?�{����i�*��cz�P�ZX���twXn(����	d5����:��?�u��a�����}w���~ZS���5?aD@�<J>��3�^B�o@�W,������/1�� 0�UM?A	�)��i�2GVQ��jߍ�Ru���dl�~z}9���<j��k]��y-KV���+v������x��XS�ī[hZ�<�I;��oF�����_�=���MP=nqiK5FT ��,���1�-���au�{lqӗ/Ln�o��T�h�S�j$�|y�6�[S�xX��vz���դ�SD�<����P�v$�b�-��ں 5Ybb.��6�����lf]P��,8�x����c�
&("��M��"vF���2�O�X�w��I&�wv&�6��˨��_b�*Gkg)�\a�{�}�B7ې�`���ৣJ��$���x��Zvl�A>����h.7X���@�O,����o���s���(���M,d;��E��d_�U��'!��<�
���6y�I1N��º����19
�<�8�����'����&��V��g$E��@Q���}י�wG�&5�i��jd�1A�OA:�`��[��e?�yn��D�0x�����n��&�ZO�W[���a3��C�=���&�y��Fˈ�w�6,f�,j�!"��.գK[_{V�msR��S�U]�:�A�%�,#�!j��	��ڑf�Z��2 p��4G����>���"{=��H_pqý&l��*&��-h/��gd,O�w���+��e��ly[; ~�����S�H�Q@��seD�t3�V\,�ͭ��m?��n-�H��ʌ�}y�@\7
2��� gl��Y��9�)Lx�rĺ^��c�{%c�������C����jr���p�j�֥����ɡם�,���+��w]|�i�?��j�9� eo��m:�A�=�U��	����߯pH�1@�]jg���A������W����VP�ٟ� \{��%�=��u|�XV��8�18qo��s'Ywu�Qk��H����.$��lX��c*�l�ᴏ�&�ȍ
'�t������Y~Y��������6O�D�:5Ǟ�✁c����*�#�>�V���N��xV��?�pܬ���>��B}<bC��$�F�ʁ�?��Q�ʽ�[N�4�:w����>��B���f����9G8�OqP{{؈�@D�F�UR헻Wʀ~Ul�Dr7���F���9�$��0��#�%��nnm���b؎L@���$�(���5{�Y�������$�66=��]�t2��7��q�������?>櫋�R��a� �f�|#hs���N�o?�Y�sc�\XaN�-ϰ�t8d�����^�%nP�d138�W�HLcp 4�@�ۋS�qC{��/���k��V)��ڦ�� �E�ъg\j�j&�T\D<!��oc6T���@&j�q
�d���nD<�OeUƈ�K��?��������X+�p�Z�i�Im�I���͢�њM�u����K��%�&r�Ŕ����E��i!��x$����u�<���gzP�U��mO�
j���[�E^C�C򽭫�Yd� ~�G��+9hV>57��n3�����G�G6��z�A�W�0�e���۟{��~ǧ�uRdx�������M}Cle����έj2}�����q�T�'��νI"L5AA�ouҸe���X*���N.Y�ypBj����2��GG���mΉN���/z����@n���T7� ���1Ԫ��4�*
p�Ch&�>!��42�����J�6\�����Cw�{ּ�hS�/o"#�/V$Nڼ%�wJ7+������E�3� �~N��WwW�WVR{}�&PX#��'�q��b���T��,�V���U�4���M�xx�JF^�nb�t��=��=KĊ������r�L��oh���O�c���m���u�D�<�I~�$����t3�����p��/$	�vʜ<ƈV{���~7:V ]hP�Ԩ�`VL+9g��.5���/����u�ϥ	����E@;F�#�0��}�w;- 4F���KX֏O��B�fJn�m�ae�şO�ȍ��l_-��\o�J+�n��n{zܑ�k�n��#�W��H��1��:�?���"Z_ͻn�����P �zo�|W�Ŕ��ł�e~Y��@NKkx�]�S4<y��p��X�OA�w^}��U %"h���) �cCJ�uk�˩m��0[��y:B���B�E��ͨ��o�qDl�e�������$�A��3Ka�O�Ƅy��?7����A��7�P>����b�ŁW&W�0�ߘ�犬�h:��]��
�]C<��R��:�ܛ��<��Ϝ|�$�KE,`7��N��/:��#� j���j:zo
4�t�~�˽����JX:3��o)ڇ0��coO�����nɮ������+&�j:6"-�M=o*�LJ"T����f�U̍r�ޕ��(��,�A(P�-�#/L���|t��)�"6`_)p�^����)p�fj,��S�N�^�EI�ۇTq��CʂG!D��l�۔�Zy�˂���#�`m��"�S��IcI�k`EHJ��̓��=�����,��Z��9<�t��`��,�^6��)3(��������	��l5j��2y�A_̓T��K���&»�:�T��t!Wŏj�{�e�A�#Z����v�(;mE��sR�C��F�>��oK=���AH���Fv7��@]���;��o&cubO��6fEA�/�����*����$�yEY��uj�cɇ��!�"��"�+��{�A'x�eY�Y�3��#���U3w�L}���엙���Y��ԊK�N���m��>�?W�TBK��7{��jiiB>%�>�_��;Cs3c������G�ʞU`(cO��;�:tK+Ti�/�ϖ{�<��r�m��[�d����b�YL�����A�uw�֮H�����rbrR�K�\?��ca��3�B����o�Nzs���߾@�i>P���>w*@t@�#�Z#۔�����SҰ���R�_���U¯�vE:��p���Xb�ߥV{6@:�g���i����fn�m�j��XG�r7v���թ�O��5��9&��]�	
�2s�"���<�����Du���
���t��5�|;��OFŮ�/Z�ĴpD���a�{v�ݖ�L��S�	�ה�Ψb�@�K�3h���[��>FR�,�����W
�j��G{�����,\{;���拭����K�Ys��ւ����#ec�\C�Y�$`Q��4�}���KțU�ԧ�v̾<J������ZY��Ye�X�"W�.t��h_2��F�>e� ��0\�#�y�8�(��u�p8j���Ԡ�B�Xt&�EN�	z����顣b���K�s/R���u�LR��Iw9��ρ��lիt�<�J���g.:�yV�gL����'?>Uۥc��2V*���3H�7w�ʉF��e��q�z���f����^�U�28�V���J�����*��\ؘ߫��M�������$?I����U�|��d��$��⁩t����>s�����M��H�EIa������[�Oj����ZcUT2��/�l��B #�p�v�����Ȯ�.��GBq��� A&f�#�W��YS%͔Y�L�\�+p���V���(S�'�ə�a;� 
*�i��2�����_*iA	5Ŝ"�\R*/���0��s%E���q�^`��./s	^~�UGE�k�c�Yq�^���8��8Z�7/�r��i8�� �пt�{C;R��>��,ԉ��e�aWK�w1�
�۩�7�b���˝�杜��-tY)����IYj��R1A{�|w:j���b ୞>�@�%s�hݵ��-��#�M@
�6ԵL���;%���kxD��Z"Wc/��ho�V��m�x�O��F����u�V||��M_�����r�#wrC4G;�l�,!~�f\��{/Q<R�)�R s���"���G�Xd� o��x�`*�����J˃:6��u��icϿ�d>�D	T��{��{�+~�����N+�57���V��e65	�r��J?�?��;��&���"*"JU��Ҥ�h" ]@@E:�ׄ"6�7�M�t�B	��P�HBo	$��@B���=�绮��������7s�޻nc�����,z9oT��L�yZ\����/I��+�X�B�y��G+lS��
�jo�&�PV���[O۱�xM�և�W�7xtg��5�(g�=BT��ɲ�s�՛�G���C�P����/��������;]�.
�� ����qng�0ڥdɁ/(�r��|s��	��d���b%EE� ��:���{:�Z<�;hv+8���ui/�b�%6����R��Cs��OMpZ���9]��C�b�wZ.���0��S�9*��x����΢<��M�B,��*h�C߇n�+���]]�?3da*q��T��9����0���6�A���\}�P1_\�ёK����#�k���2���6J�AVU���ދ���K�\��aL`ƈ��N���s�I0]�@� ����-W��o1󟆡���H�ֽ/���97�ծ�������6pA��)�ݷߜ��u���Ǩ0��D�t�'m�bl���W'��D�W��A�����s��� �W������x��m�����nE�û����Z���,�\�?N)������rճO7�=���IBm����W#S��������]\;��OƄ�/Q�(�����%A�.���>�������wX�1�(�����P��u��Y~��&�]2��:E\Z��w\�O`���Ѯ�톊ruL����
����k�wA[���K�1K����U��x;���g�Dx�i#p�$�8c��CX��n����;&���h>����Y6l%���%[����N�~�}�a����-&���R?�v퀯��>@������yF��6-�ʢ���g0��� @���~��Z�����~?��h�2°H�2�b���I�.�x̑j�E��k%;���2�M�6.��O�W�6����|�OH.����PW�sp^,�K��b�#�&�[���v�1\��$�j����C��R$�����y��V�2��_��ji9؀��(ϴ���Φ���@�\a���R��G��\��9b�'m�2��З�}g﮾�(��?�?���;�Цf�$;� ��fc���?�d����o��̀�]	�Vʸ.f�s�iLڼo)�*���?{t�� f�*��`��Ѡ��]��X�Hu0yS�CT�Ry6�H��.�~I��.��ؓp�~������B�!����w�*��~,&J�y96 HH��ݵ����*/��&O��aY�S��O��n�02RV�,
h-_g��o(�Ze9=�hW�(�ٸ�.�Tۮ(s���ӽ~�T��u?����ix*�I�ׂ�I�������� Ne�U�Y���ʫ�Ѷ�'��}�sH�N�5����>Q��j�$��V��q�+��}��p4�T��8�xLx��6�*c{��K�RHļ�ܲޯ���X}��@�8�^2W���P[��牢���9��Ak�ǻhK�\咚Ԭ}�ǳk%E7��X>p6"��z�qgΉr������o�y���E|�8�	���e�T���s�)^������2��� ��M���w�&[�a���=ϸ�b⸷����/W��&L������Gu������s�%�M Dj1N��jNw�KZhZ�?��K�p�k�1<,��� �"��<���29�����5wG�����g�K����.��?;NL�T�&����Qk���_�iy���9�Q_o�(]��ll�����?�D`������"W�J`��Y��mG�dy��k�#���Ȩ;�>�I�91�N�E����xb����x��yoT��5^չN��|x�V�66���J���������DbT$$��).�_��[�a��~^���*�X|૘ ��ɡ]�GZ:W_�3v��z���ΜCn�t&zMHE�"~�j���a�/��zse��Z.���Jܷi����>J��z4�
��k�w$�k)
W�F��܄����o�m�o-��b���S��t���JK3W���
�z�S�W��S��a"IJ�r��+��ǒ���0� �$�m,�U�ލ�]�Ռw��[F��m�����ۛ2v�w4=�<��O�
]4���%=zF�y��-[����������#$ҫ�^h29@��=���۳7�<.�Ҍ�����(5�9��v`�zb���y����	��
�����4��fW�
4����Kxl��"]�7���+��o��9����	ĵ�Ct0��MQ
���k�沕͖y37���I�<�F��1>Cs�M���q1Q��H^6П���2E�-�8G�ef�9d���/�A�Ͻv�ہ�=gI�������t��I���?(�s�2� ���E��Z�+3�\�Ф�e�uθc�K����~���i��\|5ǎq�����_��(�R�Ka'4r�6_s<��{1*-}n_FF������7���74���	��:��iw����D��Nb�]\�����p]S�Tnpp���E���W�����ij3a�-���~�<�0�s�σ�]��ӛ6Z���W|_3p���d��{����Mjf獼����klG�%Q)�'�@����w��+��7�K��|=L�1��R��k-v�˿߯)o��i�R�������6�ˌp$h	\�=ZQ>Z�{\�ҟ>�c��E�羭�ϣ�o��bN)G/�Às�0��cD�`����V�	e!���	�ָ��2owƄ����l���O�lzDL}Q����^�
G�iq�g��
nͭ	�;�U������3�i+�� ��1�����]��p�;[�j��J��}?�	�=M�Wh��%�02��nէo�������mW��Y
h6θ�t/8�]��|�^�F�	3�<y6�{a��[�@��P�t�Ux�0eb"����'F@3i-d-���,��x���+��h(�6z
�1l+yӹRv|�U;uk?hE%JOU��*Z��V4q�h����������Ap����M髬��.h��B��&+Q�"�;Hqv�q��$[9,ؙE�������xK�5��x ����d�\M2���*�B:�'�E\��_��l��H-l������j%6��eѸ�BF��Z\2��m�f��T�<̡,�ƫ?�P���V�����Uܜ��9���c_�;�P��G+짼��*�7����5�������Dx2����J���M��.��X&�n%�Z����x�!�a
/V��}��Z�K��(~�Ь��'g9dŕ�S��� ��}�SyD,��`3>���*�YJ�DG��o-sM���p� Rn����������~n*!�[�������a�9��cZ�N������I���9f6wp�L= zr���������n�B�2�lV��	� �9��>�e6�Vo�s�߮|3���w\Xl5٭.>���B}������2y%{+����x���^��2��T��Y]���W�զ}�u��_>��oo�8�ȃ����^I��<{V��2NQ+E�6����^n;�G0%︬��ͤLߘ�e��|���R�8�?�f��C�"��sai���$�u���}8�3�˥޺��d��6�o����~�U߲M�
�O�Q�v3pu`�s���������|<+��S��L� ��w~�����jϦQ�ㅻt��)���hR�
J�Rv�å���m9-q������ԎƵ���#0b��_�
������~h4�Rvs��s�LP����!ؑs2ؾL�(^�/j5^�����|(���y�H��.:/��R�Y�|����C��~88t����&���=�ցb�����ԩRo27����mw;����fa*���~�����J(E|�Ѵ��(�����!�T=�����6f&t�����B��}�O���
�����T���!����0�po=0����J�Q��{{��^�qU��a_vn�2�(��׸�^H(��k�}���( ���Z�V:z`��Ķ8Z�Jヤ��.�9催Z��6uȴђ9W��Ϳ�=q�y��h1��U�  a���C^��z���3�PS`�]����XV�Fdid����c�b��h��S7�B��ս��T8~~?�n��!w��g���p]���D̅�6��G�!V	�����M|��,+�* �<8blsE3�م6i�2.�i^���2��ښz�sS��/.��ѽߪ؊�py��G���޼�L�x.FSj�^翑�9�^�c9VՆ���ۭy�]����|�'/����m�]���5����RN>#.��O���R�5h��J�O����9��dh����}<C�)�j���-6��Vi"?C���V?}��"
HZ�U��˅�58F#+c��Rg�9����q���,�0H�C1�t������Ʉ��h�
��'(nO�%��q�UX�����H���{����׷���Ȩ&N2��'al�X̍q��a�5���k��&1�p9m�[��ᯐ�^�����a���M��o�d��`�s$�����u�ߓV+��,��~XJj^�/��K��=��s�ϝ�Wg�,����C�%F`ὭdVP*�d�+�\�����<��}c>��gyt���4�!b�ț�E]͛����'�T����Y̚;���n�p�{�F|�ɊN��wT��o/XQ�\� ���'��ɁBrݩ���9���\�����-{�:�3y�*���ĺ?�adZ�|)��Y������B+�� s-u�y4ӁaAfJ��[���A���fv�k恤)d��@Q�~"h/��[
�������[��i��y����K�%����*;?#��ݱ�'�g7�}�Ô������/�@�?=]Pc�
�MYB偃�衟0�|�q(�SFXt���)m�i�%F��^����AOi����O8����߃��	�8��$>]193��h_���B�3H|��R�~�+�=�S���̜}�:&t�+0^B޽�J�����W>B��U��.�S/��><�I�Ο��H�9=�'����h6���`��1gQ�з��J$���㙮�����N(���r�`m���ܟ��� \��q��+��2�i)L���Tj���G���RMlV���	�������`�C���aeK��;�e���:���H���E=�u?�p@�����J<"�%+���Z�1s�r5������E����iN[oؚW����<��x�L���Cq�`'W�����U��O��Q'o�T�e�f ���H;e��R��=\u�B;�	=3e~������n�"{�h{���H�����׺���Ƞ�K�X���\Y��+��q˹��ֆ�v����sQc���D5"���B@������,�2�,8kN�%��e�ty�/?/z��4z�ӛW{�0Y��031�dհ���@�1b�5��[�M�ZfN�@j1 x&1I vv��E�kq��"���j`��Ii�E�A
%xG�A���ۃ���3Iϩ�ٟ>�;Ȗ�#�wc�'��4��k�y�}񌀑�<u�aMda�LX(� �?tq���u��Ô�Gj�u2)�fW�؍i���P<�������[��l߻�D�jEy*n���3@/J��j\I�'iJ]ϓ�F��zv��M�ES�4�/X{q�]��l\SS���G�0���ź�#�>DF�J%����E�]��C���n5������i��{8H�\lu�����wE?<п�|�b<�3_�K�a^^G�������hꏶ��	.BOðO�7X?;����s��c+�h���fA����彥X����{�5��	�+��m;!�Y��3�b��W�wt���o=�՟�f�}`���x7�R��&o=0��Ԑ��[��$M ��[�9��~j��"*�D��8[�t�^�8ob��~����T�z�K������QD�N �r��ŭ�?��A�ࠛZO��]���S*W��="2�ue~��T�G5|$s���U;9k+~[���ٯ�[D� �<K�sۅB+ȋ^/q�&?g�V����2�M��R�Gc-X�<���?f1�R��Y�S��8�5��.�
	6��ˣ�E�%�����ߡ�1�w���{�_$醼�J◖�ȯI&�T��ep�Wo>[��b!�|e1y������� ��,�2n ��`oN�E��%�$/�G��G��7���:c�M	}2���v4)��髛e�@?�a��}/�=<���cؠi0T�R]���X٢��λ����ja�Hн&���Q4�����Ac�$Đ���P�.-%[W� ���=�D�M�����Zm��_3��Z������DR��Ԣ$�G�1s�����p�t���]w��~0Q:�9��8�h��e|���6Z�|1�!��wl�M����;A_Ը��[�)(|Y^~#�-��1���~g� R�V7� 0kv{��ܪ'=vzܵu�Ubmo���T~����Di��2:���i�>aԢ�$\hހ�?p��c�����n�z���A����V��a����oL�
��	�>i��:���T��7Em0`֒�kr��)u��G��z�	�L��Ӂ�f_����0E�V���X��J|5tޥ�����ܪVTXt��
{�v�SB{�O��<���C�.p�i�#�F
�[P�Y��;dE�뽱B������PN��9�����u���(A^�p���xQ@���FUB�]���6G��v����^1�&o���l��ZW���2� !�-�����0ʫ�v{G,讇��{��7�8�n�DI�^໑���aa��Ëp���|��Y+�P�8��(׵�2��3���K���3_�0�s��j�D��3Р�M���X�"݉��N���}��I�
KR{uFf��>r:�����u�_��y�����d-��[sb�ʹ��������J�^���U�,T��3k}����B0��]F�'g/���8
��j7���x<@.�v~̠ۘ�3M(F�� �Ol1�v�,o�9��NC�PT�kƮ%�
�����$��-��K���W�JI��{Ɂ��u��T�]N��z��Y����hRb�;�\ )�M*�}w��>��2� �p��]z���:��F�g�.���� �mq�?�^���8<��sŭ���p��ҁ���P�ƅ�%�����II�>����<`�E���T��O�p}/����';qǔ���1���=�2��C(����9���C�o/]je�S��V�Pcc3k��~#�x��K�*|`<>��̖-Ԟՙ��Gf#'�	L��u^��q����1e�T�D��in���2�w��w;���w025���M4����[N*�b���H���N�}���W�g6u�������i���QQq�T2y�i�����Jŏ�a�^K1�(�DH��S`8���%}�G��.7x����{��� ,�H-.V '�J�Zr"��gG���G��k���dL��f~ޓV��B�����4v�������	[�=�%�}y�hr��ً�'�=T�XB�OP��Q��3��'y^?�&�u���)r�����J/����b��v��Jj����{����Ԋ"ݭX�VL�N^�Vqsc'�� �hX�g��5���c�܎"<�
��{�}�r����v-�����\����=��^��y��t@��v�*w����/����z��76��n��ۘ��������M0~�2����t�o��͐$�}8n4yE������io���]�^$y�7���"�&��.�j�h&�OXb��Tox����3=�M�qj>#���{�M��-��7�:Ν�ww�H����ё�� {Us�Otn��ѳ��*z/C��&�Y)?���%K0@�_	Z۱���]���)���`Z��o���dQ��ƺ������'Y2��NO�<!D(($W�!,��ek�"}Yca��C\��\Dh
R#	�Zr��}�J��5���>��|���$s��j��n�z�����km}Y?0�K����sPs<JD5�d+C'�����'P��k�M��	Nl�����SEepyA��&�x��3�����|�1 �l71x�@+G�˼d@ps���zSBe���'O���QZ��MK��{�#��	/~WFg��<��H���%����T|�LU���"�5C���x���2�S���J�'�-8�W�8�6�v�>Gt]j>��PJpoB99PG��9�*.���<�V��	��@��\}ܹ�U�k��Ǜ�柙 �1+����[2������{'�Q��wʬ��/_9�M�w����?'�Ը��W_3�4�P�ٴ12��܁�e��\���`����=�0�99�4\g>�8��Q���X0���4��S�O�T�ܜ����@��.��V�H�ugV�OT�wO~�"O�X�]��P��J�"�'�C��Ŋ��/���g�I���YG�A��� 
������Q8h���S.���񷑽�Št`�v�'W��k��g�A�7���K�טҼun^�U�˞�ףּ�{��7�G�5�*�.<�>DY��Y�x��I�)�ђ��5v�~m���P>���oY���@_��;t���$Ez+'&�r��0�9L�f�@Lq�6U��V�{!��������G:ܲ�$m���w���%_4��l�8y$?B����k{n��C�+`[c�{�;+����j/u���
���TU��ɾ���W��w����"���5�}�#u.���f���cIr���g*)T\LV��ݓM-qn���j}K`vd��:;�i�N����x������65��:DWy���`�)#�^�+��:��b�N�@�r2;��%��T�����x��O2�d�����
�2A�gVG�c�h�5����� �zh�� b@Q����}��;���vO�v��4B��`�k�B�4c�i2/�FZL���,�]����m�&&�j��}}��ՍJY���B��^��0^��j��Wf��C�Pb��: ��f�
ܺ�,Q7��aC$	|��i�.������*ԩ< )�����ؒ`�X��S�껒�_~�k^7c� ���B��ٜ� ٥҇�a�4�N ��Tw�8Q�ƥ^�
~,�U������m
�f�g�%���}����g`S^Ql�F���H\���8ʹ�5��Ї#Yr�^Op�D�J�{�E�m�~<�0K���Wa6�pO���u_W�>u�x-N�r�Ӗ�NܼE��,���ߵ=ta.e�q��!�O����@�qG2�蹮RDu��A+�x��\1ƛ���g68�n�H�:\�����%��<+k��=����4-KQ�=Δ$�r�K��x�Q-y�p+(Hp��@]�eMO���Tn)"�0����z�F��7n~��ly:�H`W<������o�FE6!��M&��\���0���F:�rq�6���jRO�hl������@�k�Oٓ�R���ۙ�s�^�e��.�~(퓽R�&����p;h&��D�wU�TX0�e���.���>�[�ǳ5sw��%Ȳm.w�lFG��}nQl-���+^ס�������N��H�oj&F�yӟ�� � �S�3{��d�1���4e�����gw;Q��n5��}�!7��X2��b:(��cј�߷�[���L;:�V�a?aXx�̼a���j����������������|%�`��%���,��քK0��H�P��o�6��R�`2��A�7�����k�>��V�P�������-��-g����q��v�����4���~�i�Ⱥ,�Mp���O�� �(�8<��e�鍏gn�>B�Jt媠��*��z�vC'Z��|VJ���
��TX�CIR�i�V o1ֺ2q�i�.�Bе��������>Z�ty�H���U�|(5��pQ�L�� �SB����~���[��I�j���������"u~x��DX��@����/Z	�ө�(+��we%di�"�B�Vd 5���A���&����k|'������Q�9�5�Lf"�&�V<�&�e�b��>�]��$%&�$�!Z��^Z��/�2婝��܁��7��� �yC�G��	~�����}���鵮�V�-��^�s��Z�)~�vlx��+����x�=so��l�A-?�^�{t^	�^���~�S�^�=O48�㙯n,�ĸ}�Fa/7lkd�ǡ�������Q��#.M3��B�e�2<�T�uRW^E��FJ��7���ۦ��D��!8�Ǭ��M�i,��	:�b_��q��ͅ�%�[ߵO�L7]=VW7�h�6ϪK�فis����ָJ�����J!e:DC@������,�<բ�D��)��Fo���k��>��|+�{T��Wf|�Vv޽��d՗�(�{�����pGGRg�L���GAD��]gq�Z/�c+�Y�b��ͣ����ۀ���Wz((�2Ի�2�am��i���S/�e�$
�@�K�w35v�,hY��1Q|'v�x{�T��wPQ$[��Y�Ak��N5�&�Q�:�ׁK�O�P��D(���%�������eFK�"�7S�A�&�
?XSn@,�����e���3�[�Qysff��5�K��jg���q胜v�P�=r��_.1#�����Qҍ��2��t�Q�|�iRB��QŉLv@tB�w��_�Zm�@�'f΁����B4���SR�O畽q�i�^�yb�c�`npII���N��w�P�Pޠ~L��+��H1�E�o2'6�Wo���$�F����	�N�!� ���kg�F�η�[ ������[�2+1�#9m��K�6ǻ��6�)ms��/�t���*W�|������Jb�6��f��Qb����PN�ʸ�u��o�Q����439W�ļD@`�b��:����W��`m�V4���*+M���m|�+�y����m�pz���s��Rw����ɀ�ۖ�Kir��(�L�a�x�{�����'�j=�:%��?8�@�p�ho{�BU��yv^��弴Q�`���)��e��s�;�XmLo[�~v`����v��r�ڛ��zu�1f���y�XQP>_ao��cE��Ta'x��²��pdO���Q��%\�']h�iƪ�Qj}|cb]����} b9��'�� ��������sMTjl���H�~��С���$b�$���̱½��O=h��'�q�����^��J+,�8dڝ����K!���U�d\��#y�ˍMq��K/���y����O7�ݚ�eg���Bd�N����+ƕ��
��j��6G�)��_0��^���������pޏ���s�.Gmo��q��
�����/G���A��.�i��w*Z��k^�o�Qưf�SeY��H�A(�Ӝ�0����>mf4�ذ��.��Y�դ�e%͛���]���f��]�dc�_cM?|�~�b�2mhG�?T�^��������ˡ{�̽[t��*�Y.X�&z/&]5�~�}*��� ׎�Ï2��Uw�Ռ��i*�F��� �5s�ƍhڝ����J_'{��V,�S����<��bS�诽��F=w�b�K��ѽy~-�ڿ00���Q5'���I�g�zM�����������[OZ&%��i47H�%ϴ��-�s����,f�a��J�-���X�v��J�ϥ3�d��l��N����๗���m@��t�zG�̪�Wz�?^��<��3�o?]?�@p�vj�w��4�P��(��G�a0���[1CRe\�F���O�Q�!8ֆ�y����F�B:�#|v����е�h�E�/Rz)���m&�2��0��#��VQf�p��" �(<�(љ�X�^0/������x��E���D%k���E˘Sv�������*=IC�/��|�����s<�R@C*	�0���.�Q��jR�JS�V�o3�K�R�{0�䈡�gEw�ꇼ(΄��c���!g���1x�JAKݐLL�f-��ř��,��$@:��P0��P�U�c!�U��ʺs���K����ì��񂉟oRMc�������ݸ�r?e�gx)��\�2�� ��x|c>I/����k�l�z��p�ə���U�l�s�t�������!���s�fko�0<G��[ռ����?ϝ�*l\����Ȅ{���άɗ���H/�)ɻ�N���U�h�7�'R�*��d;�>�qA-c2�%{�H�(���U�L�oL��?F-b�l�@r̠H�D��8/%�pn7/��G>�7(���S���=���d�EC@���a�j�J�j�xW~A���b�g����b�ֱs�3i���k��1Q�%T/�m�M��j�.�vC�j���׽*����g�d�C�~y�t����P!gK	�ӗ�#���X�ʟ�u�J�1@ۺ���iJe���u��_pyo����'�&7�Z<Q�Bi���{��NYЊх_Yq�&�5�YY��x�D;:��-W*��G�R"!g��2Z�J�z7�Y]�[�|������b;��{�>�%���t+�V+���d�T���`偪��cg�+�+DP�*��8���h�7w�!	d'�"�3���+SL�V �]����A-c:�h�DmqP���@�&�mlg`�=2K�6�Js�4�䉑rN���!݃���l����NxC���6�6��=�����̼��Yy{8ƥE���o�w�U��M%m���Ɇ�8=e��w��>h5H����I�����Ҋ���
갫��gTky���\}����G6�!M������gD�P�V�{��y���������z���[�/��Y�ܨ�}�I����'��12�i�|���=�!%��Ӈ)��^�|����M�_���ɾã����e J��"�X[<�<�]{H�����,��Ї0��{��f3]�J@�!�	��ԍ�/�{�W���M|������>�ݴ� �6��X��`�&��FL�u3R��v�=B�k�S7=�4��F/��M,����ǐ'EL:�z��MY�f�n��I?uQ��*�u
�;م3�< �@�"e(<�&�/_nm	��h��=�H�0�Jn�-�:��/�`"m�	h=��y��N��tp�M"m�;:z���^MwY����d�}|���1��w�f���{�(1�ﻎ�P���L���"e1e�Ѷ��c,w�	c`�ؒ����]���'�l����s���J��=Mϕfv#�rZkwDxs�������۳���l#P�e�=�	�A\�a�HO���|Ľ�@&�>�D�E�g�7X[�z�̄���;P���Fr��ш�� }m���3���9Cj�QWʚ���֨��_��~ǷЗ� 3U7� y�s��]9�y��n�O��ma�߫RH�ڔi���o9G��W�\s��@.�U�C��&VP�/+A����LxL0�mB��Q�L���������R��KG�bF�.�΁>;�p"�PZ�T��6�1�z���b�X}v���tb�/�%b�nrO�f�;-23��5T�٧�L֗� �|U����K��ֽ����M|x^B#{~��q3�� ���z�o���5j$,�`{z�9�~*C�!\1jѫ�'�_U��!����Č�GJ�{O�,6?/����� e���*{A���{�&'��v �*�FĐǾ��m�kIᇮ�(����^�tF�\
��M)��|w� K�(?u��?+�,8G��y�ͩ6o3��R��Q�sG�s����v�@�M<��<^c�q1,%+�V���qk(����Q������>{��=�z�uOي�d1E�RUe�;���XA��V�'��o坫���?ި�|�x��%�szzP�x�����0%���4��R�y����C/��kg��K�mfm��Fw(��닜�y�mőR!����$��#�RE�%�N۩<��I&�]j��K��|��v���z9������ *���k�R��L���Tz��@��R�0���3w�����h���B�x�8��24������3k��kI&��ĳ"��,�`�.3~���T( ��Tc���hպG����/lXFe?+B)A��2�Br����e��НNݛ:~tM��ԟ��j�/~1�)Ȝ��ZC"X+���j�cZ�YҢzi�I�Xq�B.�8�6a����תԉ�V:p�7v�� �d� ���*��l�=T8���P��J�Ba�AG�`6ҙ�5�lb$%m�q�^���%�O��]����&���e�k�Kd��ݷ`v�losˬ``}�Ds���V�hDY��x�ӛ���:��}��&Iy;2��8������c�wd{c�-��:>�0����K�V��7�С�p�dqI��D�C��97�(nw�C@��S'+-V���]�t�˩'+3c�u�|e��\Jen�斉V���n��jb6���rX �T{"2۲�)�魦�\�M�0) ���7�a�Ҧ]��;x��݌pv���]��	�
Û���G��W�?�D�[Fq�ޘ"���{|8��?���y��Rƪ��Vm;>VO��2�|蹁�Ӓ�a_�LD*)-PH���y�֪�ܚ�2>w3},E���̽<�_�v8��Ӫ�^�~\�&ei�����ͳ� �x���EvD��kT��<V̅]tx�����k`��Kc�[g��ǥ��=������3Z���r�Ik�Z4�ғV瞇���ب�])e�R�a�2ؤn%vaU*,UA�۴6i�!�����J���Le��8���A&�<[4.m.;�؂���������K_s5��]��ɜ8��R�-F#�ջ�ߣZ$]��C��v�?�`��I������Ɏ�+�-�64�q���\���WL�b��M8���R��W���@�@�\���[����q�F�V���V�B�%N}C̲�ֳ����g^������^j_}�	.�"z��J]���6�\�,#�f�A��8�-��Q��¬���ew���D{�>r��.��f��t�^�f�����8���Ϋ,��@ɷV���rO�K�����v��]W�[W����hk�{g�m�������) ���a��ʬ�Z�.10��B� xM֤[�"N)�y�]?0Q;��V���@�|��,v�&��L/b��A>̚�"Ƴ2�'�Y/^k;ٔ��m�4�;c|���V��ŵ&6�]8��@3����X�^�E�w^�׏Q��f��h0|�a!E��<V���Q����P5;B��mi�V#�ƌ ��E.��E�V����)I�QW䚄\(@��o]\�rB�5m�}ޛ���ew��o��e �������$:^�7\��,�˂�7��N��E�ߚʝ�,wMϞ�:#����4,��^'�U=$�⥔���4����j���㛯��ޛ��9���U�ڥ�J]h%-��3����mI�]@G���|������@,�{zY�<�3i�<RV*�LC�#e$.���Md����Aty�����vL����8(7���������3��W����&�zG'jc�D��j`�_X>M���spG���]=�C��tq���K.�9zyP-�;�k���6Ri/�{�0ikۡ�Q�NBUJAԒ��-�������m"����!�3�":�?=#j'�QT�D���?��3᥺���	##�S��T�	K>.�^���	{g�#+*� �{���ο��x�<��.6e�%wP_/.�w�vV�5�1C��mR���e�;������&F*���J�a$$)E�����a�j�t����|?���2����n��;Cdw���a<pu����p}����b�ۘ�e�ޤw֏r�ٚ|:�r���c?Q�������v&ƣ�8���MA�����k�I��� ��C��K�5MZ����MH-"�g�v�IK��3�f�$w�����Y'�x�g���!�'P�����Ҩ���V�wr�e�������׸��Nf�B���.�h�8��_�'���^1k)�J�s:_�������T;,�RH����X]��*�5�q�1 ���d���pM��#iJfQ�Ff4�Ff�+U0/�=8kȂK1��Z+�����̋�YP���%$ߞbU����{��B��+[�~��`l��G[��؆�� �(<{q�mʡ7�����ߕ.�x!TLq:�M�+�ʯ��%����wt":���Z����T*����]�k��N��Lu0�f�:�o9��@]�������Ύ�3�i��k�I9�l{����q�,w{򰀫[�{xf��'-*9WChU�ڌ���s�����S#Y|F8��n�|V��Y,,P��+��+�u��[�n�Q�V��E����X�T�kT0�~��r��TRE��2рI/���
>��V����g���鯧�$���X9.i/�[ۻG�(oŊ
�%��ae]�� ���;�&āD��'Dn�#3�Vd�˼�`h�ޛT��)/��g�}�M�r�*x��"�yr�0<�q��HM���E���=�`n�����52���r���~�����+w�AU#O��5s��Bx#&H���c�i}���
�8�����f+ii����Ⱥw�ii�w?�O�R�%|)a�/±{RuE�|��g�ħoE��?����D�ǾT�`6A�:+�uS)��cb�Z�0��W���B0��y�'F�'�j�{��������$t]�p�]v��B��n�Hi���M�පF�^�y�6j�c\Ԉl�IY)\��L�@J��Ş��l�/���8<��������n��g�D�m���-���ܴ/�Ȗ�U�
���X�L1��Y�Տm�K�u-��iMG�����ƿ<Y.����d���c�'Y8�����?����[k-��d��C���s��.%T�R��MW�|�\���xE�n ��N��`�.�Uo�������8,�!@�IO�xF�W�ش!������P~o�Z�X*��"{����,	�CH�ƾ����}˞}'��%��ub�!�c�a��}>���iy�^�?f�s�s]�y_��9�}��{�'�a9�"a�m9R�P��;����q_m'=�H�3U���!�^Jc���L��Qwm����M$d�6OrJ�n�w����h�^��߶�o���^��J{�"���U���C풼���]@����r05��"�	3�^��ަ<?w�ϸ-�����Q�����8��1�ŵ)�#Ϻxu��'�{�5�۳��!�� n����x��E���q-qWe�$ɼ��)��|9��!hXЏ�)?C��� ��K{�_+]����,x�H��R��\Tm�)<�Ձ��f
8��!����й�T��$�ηM&�g�:���]�:��),2�(��4�(�<���l�0a/��ggNY��ԓ�Z 3�KdDAC 1GĝR�%y�a3��.��0�FK®�rzRJ%�*��6��K:��r2���r���JԊ����T[�hїuѣ��X�SE7�-����^x_�6���U.s!����οm(O2�xy�2�-jm�9���(�jи�ղN룊$�����g��J�(`�o3E�=8���y���6����z6�4l�;��� s��2�?��d)�s����.�~�X��8�dz�&&�&��}dȀ���p���ހ�����8 <U�\Y\w�2.���KZ%�9���zT o}����2Fk�ǨF��1�OP���m*��ZE���������8"4}˼�$������zTb~;5U;��n	�-\E��.��D�p�ɢq�����~��Р9���%^����m.���*e=u3�"7��;n���/�6:���*�S�Ŏ�&�}�|��Kjh�p�1����]+B*%axݛ����[��k$4[ك�PN��g����־W��69/�%\�k�(y��&���2]��LY�}ѓ���1���/��"�<���sz��ܓP-	���9��g`⚽�����xiX/J�k~{����Cy�;pV^j�n�M"���#�j��-�`�)�dk�"�=�Q��TZ7UxG��'Jb�!@~�Z0�[j���s.���m�s��^L���Gއ�����j�&�u	="U�7��;�����J�;a|f�7�� ��f��P�ur������f"��9�;"L�_R�봥>t���)
(����0~��?���<�a��X�Y�_X辴��Q�{��W���?Xy�QO˲8lil8���E[��VD�Y���I��5[n�d�|�Z�v"F��,�CV@C�=�3�Э����7$b��uɫ/C}N�c#�ɱU����a�b/���Y���7�F��I��Fe�|������Zo�^)�����nʁ��\�2�ʻ���z5bF�Fp�u�*��`���u��Jy�۟�zܣLK�_��T�k	陔LW�SٳN�ɧ��Pm�%h���Cw	9���Hؠz3^;%�}<��s?l�3��>�W�7�[�[��������ݖ�ӫ����먔*�:�zh�q��P~���(ȞM#G��"�����k�u����[�d����5�/����œ�ip���?F����*G
'��r�x+|�f>?L��2�i��g��:���\g/�8�a�d~Y�8�g�Y龙[䀾�X��5;�u���O3��O����"Tȭ������̪�ڦ�5���g]��㘯�0֛qd|��� �=�y�s ���D>���Z�mH�6��\�ɻk����J�F�F9�e������U�Y'|{�B�2OSff���o�tE �c�j���j:x�";��������֙��r����!oH��*3så�I,�xb5���1�"�![�z�9���`�n+�o�*{sj���iy�u[���,���G��<�'�R2�V?�y���>�to����XH��OXG0����e�P�؟�&%ת�Ld{�z24�(�#�9��l%�'��@g��ո *��ɴR�$��k�l����Zp����n_�FV3���T��KH��G/�G�!�C������@�H�8�D5��Η�y����2��A�Eԑ:�����D����֠��a����T�7�$?��1H>&T_j���10 �w���h��Sa7�yp��T{]G\��I����"��x�/�e� �~"^��x��S�u(L59�?{sg��^���ݝr�I"��8D� �$��������j�P�ɀ�?حO����~鯙�*zW�<z)1�.����5�s��'����ca1��*O\+�U &��U�����)/�o���O�Ǔ&���C��`�7YN�⼂�`Ҝ$�"*SG���h�V��4Z���H����ST@�!�r%<�$+=
�_,�V�B�g�,"c��E��� �0��1���	�r�g�?�۸|b�%B{�|�JdX*��C�/����*a:�scƞ�0���������UQt4�㊗�?<Y�T�8���� ��{�?B�M��7�C!��W�DYȫZ��
��1�͜F����/a_�$���b���k]+$܌��O���ۗ��I��d�X�o�H	�`y6�|/������[����9e�K/qCҍ�b�ţY�&CK(�Y�m�پ�ɢ��gV�DDr���O���Z��o�d��3�61�}��HP�k�`�7���pN%��5���Nk��N͆������$dC�S-Ue=Ge��k���G��l�S��?�<�<X�_���c+;����gk��~z\�D;�(��Q�|����똅ϟڑ���	d!�6�	�XZ1\����i$!�8����ǎ��F������=��?�4k�\�������L_�2�y�����Z�]���tUv}��eC�%}-:)"�}Hz�QË�A
�^��iWnU�~�I�2:ʤ�tF�/�jUo識t7�I�v��SG *=�z�co,z��F��T�R!<����D��W�>\�������J��Dֺ9�W˞{�H!��"aa��Ź�)����ޮ:h�^4 &���u)�s[�Nh�)�_ ����d�@󘪭��C8���ͮ�j�D�;}LΨ��p:�D�Uj^�O�+%�Tҳ�x��{�uϓ�)�멡��b�g�4�4��O�wm�(&�b�jq��:�5m�@�,2)W�]�S������r@�'I�8l؞.WU2PϾ�;IoN_��^6X6��ݧKb�@{c~n'͇,>w�X�[�)=�������;zz��M�Z�P��s�{V�;Z=�X��3��X�.��\�Z%���DW�X�z������'����J��$��:.���ݦ�כ�d��{�S�M�e�*U��?���r��@�[����������
a'.�2�K�O� �JW5�y5A�GD�+¨�*��$��J�Tm9 O�O���ޟ�[;��H̹���s���1ڐ"�&�ݝI��C�wk�ߏ��6�˿�k�d�Ni:A6�����n�)扴�s�[c:�`+��;�1(c�����"2ȹ0Ҵ���I{'奥5&��l�7˵>ݬ,�}�oZ��\Ԗ��qQt@�
�ϡ8�"�Gw���,6�6f�Ѫ���_��x0o��D�cgC�������YG15���k$��
K��r���8��'4H��(���z���d��mzL�:��<��=\bf5󭦆���ؤ�z���0�ҠN&W��!L!����;�x����}�F;�ηl�ߙWx�f���d`SJ���w���|����F�钡s�Ҡ�I�����^r�!�S�\�:;�@P����B��N?8G�������Hm�;��lP�N���>���f��k��OÐA�hD[�g�f�����e��)��Q���B�<6�ĄI7��P]���y}����8�K���
_t4�c�����=��*}alqL��K�>�B�oM��m���'G�A������dD��vW����t&a|��"T�o�����߳��aV@j�*�w��0C#8\f��|,��U��u����ȯ��`&��ˍ
�0�K9�X�d����xY���N��!���
�of��&�լÊdr��fd�5��%Z�}	;�}�&����zߵ��R��r���-�q�/U� �ŻŇ�,6A��=m�\߉<-5��dWQ�^�(�+��h3��c�����/��f��wvc�U%8<$��Y> �M����>��vw��
�6��C}YeI���]��}!�,Y�����y��T��Xb�'��z|��z��G���}�!x�$����l��n�+�y����n�*�'vjx���$�x��\��L<Zl�������m:�qIw'6`�q�j:[y�O^� -����z����mi��ɷѼ�����gY$ �����9�?��zd�>�$���Eǲ�_�Yr�Qغ���8�+�p�tCq�>���"ɬ9Pz�)��c����;r6�l5��wҜ5�E�a�u8t����� \�Q���'^��JCwC(�TN�)�8r�(c�E3�����OX��j�����[	�o �D �\i�����W�n�P)MȠ�%�n�&���BO/��Z�׽2͛}j��KN?\�����pG�CѤ��
w��0�3�R
���^��>�>]ug
.毖���*!���"C�!���b�25�:V ԋP�*W�vv.�Lt�$ۣ
�	p�+&�?Z�\�6�@��L,�%A�1�/ �%r6o	v����`�#V����ӭ�w��CH�ia��B�#�B��屡֝oNzPGA����y\��[dā"�o�=��8你j���Ͼ6'��ilm�8��QI���ۼq�vP�������8yO��� �`��J��%m��,�!D���3T�Ν�7;��3$�⊝"z�F����]�=���9dE�/-�/�F֔$������8��r�A����/y�^)SE��N���-�Pe���;�7V�?7e�߱C� _5������_6�R��Lk�uX?pXA/���ihn��M���h�'��	zX��ù�0��i:�q�Գ�H�3������×>r�yRn],	:��Zq��rLC������h6vQ�;]��r�[{a�'�˺�􈏎�;ZWI��%F_��a������c՜����2noK�N`8XB�m�$rc���a�,lr�p%�T����2�JX:G��n[�〤z��%��U�q�t��A���/�Ug	S��K����g���c+L�r���!Hf	���U'��k����{�D.Q�)��*�Lc�����I)�+�ŘQ���%XU��ݍK�!I�������ɔ�SN��!{5U>@Lm#l �׸�;��Y���=��q���7�_�ˣ��l�e�xRZY�{�c~M�(��7-���O�%X��)[�&P���{���j=q$��
9IO�'�A������G�?�^�
�4G�S���'���A��B�5o���V���#��!I����A�;�wR���ud�xҋ5�^9��A��H�T�]��=#)��A��'ft�7FI$�uӲ^ي�-�TX$��gN�3U�������s����jZ�N&wӞm���^,��� �B��g�ψ�\���++"23���0��4��Vng����V��64��_��"��H�@;Kɵ��A��3��,?�aT1C�<x8c���ҹ'���R[���\w�E�+�v�G�4����0s�r7Ο�]fv�ʡ\|y�}�pXkcL�qQ��ՔWmɰ$��I1�����P�cf��'m^�t�B�=�3�	���m����"3���vq*V�L3�l���D��.[�r1+�)f5�p��VF���@�鶁b��m�~�\��>�������5��҃u��R;����,�} W�����Y ��d�X��1���ڈ<l����*��DS����SF�ߜ��sn�?��0�(y�s~�����3� ���iYt�����������,츔Y������F�;�c�a�׉3��ٙ
��ܯ#39�cu}v[�b����öZ=�\b.{���кk���h�43���h&�_�@}?����q��!u�j~t>%�7U���d^�9+db7���HG���q6&�%$ɏ���9S�ɿ����6��hש�%Sf��G,���6�p�`.��S��3�ajb�m���o���JK=��ɟ��`�r�I�1L�y�,�LH�]B����NM��6s��o�aUv)C���g���I���E��`�窖�3ś����c�V�f�zJ2S��ƚ�O*{
����n�n2��<�Tz�� -�c�K�rkk��%_-��������>hn�sE����v��v��@��#�^|�E�s��n��J����}����[��Fu�Ź��[��G0�cU�چ�Y_��p*�����W4�vn�#��s�����_��v��í���9` �� ։ˈ�8�+�=ѱզ�kYo=e!��1{-�Gw�ߒp���|�y�uJV�	r�|��$���z�e����n�_�����������r�9�RM���HQ�~�{�s1��k�+���� 3H���x�_$
�E'TScK��!��^�Ӆ�N{���O��ϼpFԟ[�"����z�u���G�5Y9*��{3���t���w<g���6��#*�P	��2Mi�|"��N@9uw��V��\ٯ��H���Ӌ&^]����B�RQ���UWY�s�g�hkh�դn'�/���	2�n�
��2B��5���s�P�Sr��Єo�U`DV%x�d�DA�~܎����@S�A�m����M��A����~%��[���i�(���C�����*��6R��o�=
��b'���������0;7�Ǵd�2� |7<�3��s�M�ѕ���"]SG[4���/�:1����܉�$���LNP=@^�a��}<��X����X���kh^P60�2 ����%��]����A�5GϿ��s8������=y�*�/.N ��z�'�Lٍk����wa�ƅh��\����ҫ���;�ƞ�1��Ӷ|��=\%ص��k�m�u:����>�@W��f�� �����������7&����>J�㊻��b�ߢ����4�޶s�*bw�qr�哊��04;{F�T�~���/D��9_��ٿĞu�ѓ�����[�7�i�(�A�a������35�g���j�hZ���W�>�y�Co��ޚ�~q��_4�����v��,���Ѱjj�_Y���K��墰�?j��8l�겣T���\��A�����F�����6v�,"�osd��_%���ߟI��my����E�S�������dl�3!�"ؕ�n�	�Р��������ח�b��[�'�m��yW����m7f��`�?R�PV��Q�悧}���2�w!H��	g�EB\qs��,B�����!�U "h/�`�ܖ?��4�R�:&����\�R����_Օ�}��3Cxqd\wRh�r���^S��m7w������2fB��� �.��1 ��P��B���W����$g���斏��3L�o#�!��ȹ�FpS^�妴�v��՝e��;�ffڕ�T�}�7�B��K�<���unN/R���ë����5�+ (�BM܊���?���7��?����)�A�������_w�Φ�5�K9��x�U&v��K�Y kr�a�$*��UϠ3���{�ĉ����.3�4��SR&ھ�4:D�ov(j_�k��[1����Z��B�-&��.�Ðw��Y��z��V�6�̞o#v���U�[�;�앉�.��%��V��D�&����\��(���j�Y~��/���kˠ�z��a��K�F �^�$K��á���3N)�G
��V�d8�uZ�ؖў�Jy���I���!a9F*��m#���!�����]j~�e��n���ʁ�)���Ȼ��F�x]ժ�H}<�����d)��kӁ*ݾ4Ht�pn�+z�`�k?� �:���g�v}�$N���NFϤ���=��&��f�������}����u0V/�w�����i��o� |��j���!�c�-���8䞢����]L��[L�ze����M�ON�f7�DEr]������A^x�b'�H~=w���ZRĤ���z1��ŵ�fn���qf:]˶T�� �����!�$�3	�3�Z��e�u/w�~��]�3�D~�QV��H&������T�l���ڷ��h����=~ձ��Xre �W��Q�a�ǵ��=�M��J0L������"ߺ$4[������Obw$ �Ƥ��Uf�a�Wֺ9����k=���?�wٱ�Q�[����[�|v����.H����R"���W8<��l]�3��~��hh��щ�ڇ�86L�>�Zj��G�r�Y��crQRd�=枏sQ7ϩ��N��ƿj��/��]�%�ǎ9H�*���$^�ջ��s�ǘ4pŉy��mlM��oh��ߢ�tf���љV$�Ez:E#�ohXp�`����ﮉֈ]��K��JJ;x<�������-|`o�]CZF]٪�0_�w�w�,Y`�^�^��&�hf�&�L����6e:��F����GcW�4�� ���(G䚪W��?{��>���n�[��ajz3���/e���,7QghE�ʖ,�����P�^��s�����/�Į����a����T�U��3a:7
�Ǆܸ��F�	��$3�ի
���X� ���k=�{%{z���BXm��i^8h���n&}R�7c�B�v��r�W&�}�+��	4�$
�7���|��Rs�o��ќ�:���z�Q�����ᷣ�P7h=��q��:���ϲ�<r�Qr�&��'�r��nUv����Qz�\I���'��A^kk���m^!}U�=D� �&?�7�a>oe��P�~��W�5�Z������S�p.3�q���K�E�"���z�.q֥�R)��X�K��b����Z���0D��p{��07ە�a])[��+5�TjxJJ��X�������[	t8BUA�8V!���^���;� Lī�v��ܳ����^���;;�o�u}�����e���h� K��h���T��*��)C_K�)"8.~7G$$��9z��+�V3��3Ӻ�\'�vC�IC�;�}O ��P��:����o������N�$�v��:d��È����U2#Fb��ʲ[S���~���n�(��έ�������2[�
)63�E��'.^+2��_�=C�~qm1��X�:낟���53��C����F�?��G�c@�[J(	�h��l���JU�8����y�^�nA� �Q|IU}�z�<Ӆ�yb��(ns1qr��������'�r��"6?N/r�O��P0#2�Y�M�O�����i�
AC�%m8�xXBxx�vh��;R��k��?��rdD���~���},��q��(�}���_�Ow�E�>(��8B
���/	�/�>a��B��˼W�gPk�Oy3�/�f�vqŞ�����=�#a��_�X�����j�[�����K�}3���c����o�T�'��l�T�I�욄K�8t5l��`9@��{SKico��ߟ���\���z��^�V�}Ҡ�Į��B{�q���=4�>���CgG�Ç��>ճ6?��cY8�8���U���/Ͼ���� Ll��"9ެ�6�����<�HrVw�Lx;�?]-p�b�
�R���j� WRWU8f݄|�}/��؃����O�z|򤾻�����L�7r�N}�7/J�Y
0\������¸��t�ϔb�o�/uU�X^�~"�˧/��؆f�)��'g� �D 1�͓��V��[}�IE^�j���jn�~{��a�h{<K�m�(��m�i����]�~�.��N!j#���'�B`׬��1b`�r�p�>%C��ޗ�Ւ 窨����]α���"�h����d��ػ��[Ţ���:�E;�,�=?���lӍpY�~w';	Q^X��2:(��|JE���O��83	��
+a?��0�����Pg�xu��
�m�©w�A)�iw��P���c0!�����v+�#�~׍�+�h��� �
D�ɓ�Age��=6�g]
��t��d������*�[E.u"M����urŦ�����-����
�#|�d�o��e�Gmu��r�55
 dL����B8���pc�₰�"����#�c��W�h3�je��\�y���7�s_�+%�=ӛjU^�X��b^$�1^!M�q�u�.E��4Cy�g�$�z#�Q�+ƃ��K�ki����	TT��ih�;�Q�0�a�x[e?ƾ)Ǜ ѽ�r��U�m��O�%�9r{I��:���%HS�?�VQ?�>�����_tw�|o�8>OGƴ��9�e��{඿����@Au���f	x�	�^=��,M�ز��б�*�F���aB��K�S��$��"�5��wrD�K��Jm_��7�����{�cK������ ��?Ti=o�8��Ye� ��{:���m���hM�\o�~���t�2��Q�v�@u)Oee|emw޺���#wy��uϘ�D�H	Z近�^][{#� ���"ĝ�O �:Rz��i!!Y�����*7>����*�w|?��O���D6tU
��,.�<j9��e�L���I�ǉ�]�ϥ�:��'MV�R��9m�"��_b�T���$"��կq�J�"h!]-{aɕ�ė	6�a��[��h�sԦ5�)����T��I��N5�e�a��m��Z��8�=͖MF\='UZ����1�0�C�EWԥ��P8`�rP��Ho\�Q�Y�# ��M����TkmSS,C�bF���^��B���
� �TA����= )к�d�]�!����� �>!a�\�����@ev���,30�EN�S�8��M@��ܤ{���7W��W�c_EF�V�vz6!�>��:?��G 3~Ӑ�pm�,��m��b�7��k�V���L!��0�c��ۏ���u�߆��Q�/��ˍ��v�A�B[#��Ml�F��� =4/�N�?w�_���N�Y�{ �+�Hj�N�ރ���^+$�hUɹ�C�����}����[`�߸���+�w7+�� �5���p��F��^��5�a����xx�r۫�T��p�N!�v�=1���e��#���o���+����Jwqձ'���6E�-G��R���RX"F/�W �=�qt{�@k4�T-��t��,w���ɮ�!��k��DGi	�����!?NpW�;�~�~$:�ᴗ�&�&��v�ʑ�	�'" 3�2N>3��1),4p��k������=}!�W��c��1~?YX��Qg��VG��d?�<�>� �>Z|��1'��T�1����d�!��L�=�����"��
��!	�ʂ����{k��u���փ,��$�+)��+�Ȓ3� 4�)�o��p|`U��s�n=�>|�xc�߯
�W���d��Z`X	�U(�&kD7g̺ `&��%7���e���E;4u��7o�L�R�����{�`��;��|y����Ω����-���~����Ʌw�a2S�}����N����|R���^� m=�n�Z�,VV!��%	��!��m�|�En7
��v�gǛ6�SM�ߛ���p�8����|����xgdf&�`�[��w#��^E]ٯ_O`����ݺ�pt��� �J!�C��9��Nn&���`��m��@g8~`ӏP�7	Ɖ���Y�-/�<O��G���������GI��Ԍ�Z5�7O���}sL _a���y��?����Y� F��Ef�0p�^��@F�y�DC�n�,g��>z�w��w�����i��4�P
�P\��X����b��t�B�1`^?���S/���)����?�o�Q²Lշ�����V�_�bb6G�z��>��<S'j��~U�3x&?��rJ�8SH�Dz�5�Xroقg�5,����!��9� �(��V�^6/��\��h>̷���ۆ_X�':P�#o��S0:�[dg�(�����Zё��`�2Z��.��[M�eF�_r`Ō�η�R|�wa0�#r��ߊ,g�2���4��U�Pt>#�mƛ�+��/��ß_э�u�2-iܘ�1�~��{DLQUB�;�������>���O`,X�� g%o;�(k�u����G��Q.�1�٩�e@�ސ��Xv E89Q��ԅ́sQ�u��y:'\"���ť8\A�C��5�sOڑ{�c&�I��#���*W���8[�d7�Ւ��аo���9<`O��0[����uU� 5ƽ5h��V̫�7�Z�z�Q6l��+'��g���o'��b��?�m|�#��|?W��>�����3c2q�OF�k����ɗ�8���L�3�R��VS�>T)� [�ii��2���S�����"�y�B��_,�����Ac�}Y�����d)��-�oD�G8�I��ޞecJ/�'�K٥�X|���]:���E��}����׊��)�%qx�%�����i>vaKk��d��R���bg�ƚ��g٭ ���dЫ�yE�]*�A^Hu���_v�6�^�+�#2�w��� 5!q��측�ٵcVab��\��N��lo@/�\��/2��W�ݟj̞���g쓐�]�?ބ ��U�M�yē�>�>g��ӗry�X��/�vG۞�\P��SD�`����+_�6Qm��]©�
t���T�Xx�����ؙ���L굋�l���>���IW�z8�x�Ճ���i�v��������h@�^�ȉ��[ ���Ou�S��(E8i�9(n4| �<�*vM:)�ܨq�g��WR�8rG]A�C�ݕ̖q��y �&)4!ؔ=L�f�x�����������V�W�@�U��j�.U|_Z,��QbcEf�E~!Je�ށ�u����|�c<��_�t�o�\7C},��wBoS���͡��_�8J%fm�$�/^g1,:k{%;�<�r��q�B����8�cU��_p0<��.��0O����O�'N#�S�@,o��H=Z� pB2�Ln Y�6<c�7�%MA:j�) 6ꏶ}�	�	�����]S�����z����-u���:_��,T��t ��P�u;6������GD�rG��$�8,���xj��+�ng����\��y��O��A��^i�W)~�*$�L#�@����p��vcv�mSNy.�H��;�U#���ܢ"c�8c�5�C��;�% :JV�Msy��O�6��"�`�%�����u���kv�%5H� ]8�`��9:42QD����*��O�����>�A]�\K�1�[��|������O�'��ǕG�W/:�u�Z8\�y�L��[ۼ��Y���/M
P^\���b�jw#a[��@��> �[�j�!�_ ��8��= r�6+1���vgCw5,�v�*6'��۶h]0��25�Illh�[�y�*����joE��/��lNq������br4�����JP2����˪Ff��������5�� �� ը���b:����w !8UiՓϯG]�g��Qw�Hӈ�a�.J�#�=YMڼ��E2��S�	[Q�fW3D�W_��P��	��@�paI��gT��O�$�g���f�}�Jw|��Ŧgq���c>����l�����+%p�*Z�����ZZ�ُ�G�%�sNׯm��\]0�{L�L�� �0��S����w���A���L�"��W��?�Yļa����θW��8�Ƭ�~���b��E�8#�ȧy�������>�ys	YO�LK�D�lW�`��]�罢��b�D9򊇉��No�����#�ڝ�c�`�X�����6�\��ّ��Bv���ɤ{ȑ��[�����C�u��CE5������㳹���V�[7�;+�����fϕ25)	�}��K���^�΋�]$��")t���X~h��  {r{�,�bC�
sz?�"�pc.l�!7�޾qu)�?e��T�܇!Ȟ�^j�d��Jc��:g���6m����ƙ��L�J�������,�4�b�_��Xi������'4^��K�iloYY0��}�?�^�-3X����C;�Q�b�v$=��	�j����{��bfVV�6��5����,��@<�(�%Ls������� ��W�` �����O�$9�׏xV�5� �������I���9��?���.�;��m`���D�wg��3J�~��IQPg�<���b`�p	����Y�8�C�����3�%qH�	�"�p�I�UG*k,5����/��}����ެ�q��`XYl���@ |���dc����#RF�7|�V&�������f�^R?Ըo
*���ظogH>s "�zX�I��� �-i�D"TޮQ�?�n9a�˗K\mƳ־�^���j�z�uY��c����S�>�Zf�����~�-�L��v�������P����!'	4�M]\�y�g��Z2੣�V<�n�~>��z!�V�-�V�bWb����wJ
�{�q;m��-w��7j�ipɞ�uo+��"�Ӯ/>�N�}��R)g����G�_l.�T�VKq�������W_�H ��t:6.��1C.N�[&%��-̍C//ns�x�xY�- �6V3}���/뛯���yo	�~�ɑ����#�S/�[��|bb��O��ǎ��C7v�x��M�+��4ze�$RߝrT�������>�
}r����N�^�dwTGӦ�
�ގ���Y[�/�u�ǟ���i.�q}�O��B�ѧ���� �������.)�&	���G�(��|H1$Ma�mD�	������F���z � �H�՞��o ��{+;��ʙ��{X�(Vr!���phwx�r�u�=�vT��X �y���άĤ0G�ON�&8!/%'I�������`Wd�����p dǿ��Փ�0�=@+��.���H$�@�LMkQ�?�k���"�6��>�)'�E��=�v�2�R`j�����VI�I�������oV�S��O֩F�"�L�i���/0�Otҹ�Z���+����(Ŗ���X�����1�������^���:�˥���v�&�Ҹ3��E���=ϩMw�>c�{�q��~��^Nθ#7�^�r�j~��)h�]=	��r����W���/>�G�.�7�`i��>���w�]~�o-\�6]����L��1�z=��u�T�gd)�`�s��n��S_��i0����i<�±�P�����F< =��\����/��we�}�s��!��P��/�a'��.��D<��5��آu�Î^���������QEU5��QX#ԟ�G_c@`ph�V��Y���׉��ܽV����Iƚ�����v��js$��禇G��ָ���hbr���1Ru�1-&�=@�\���x����y�UVŅq��>L;w�'��5.�7F���V�5.J���yI�#7�!�/������e㓿<�pW0Q�����7Ѱ�Y�J��S���A U���0��"eJ��}�~�Ү�z7���É�j�'A4�	v-+S��R���4,I���+?0_9 ��]k[�G�jVAW6en ���3��o�"�D���X߾��=1HK~"ԜE�����لIp�F�?�3�[yV�������N����4*e3��CZ�w�=�t��	��g�ф�l�����-�Dp�æh3�ed�{F�@�S�~�o��yfvLЃ��KNXH��W����a'��IL=Aq�C�,Mm��>��"��G>�"��+�+(���I�.E��4�̮м���K�>mGn�
R�r�q�!�i"� �tt	N!�z�Sd��f@���9<��[m�Q�D���p��?I�iH��D��p��1/���da�Ǳ������mz�8��'{�%Xuq���]�?BT]�J��ݥ�����"+_>��_�����P�N�`�o�%�pCɖJ\�N��9GZr��#A�}3N_��SD�u���j�D���u:����)&�N�j�t!݃����Z>O�+���^�����_��J/��cڢv�*�>�c\f�=6��ж������v�(�7v{�v���{�)�ԡ��/�*[U=ās%��XУ���ئ=Q�Q�[����_ކ��r5���U��5y�Ƀ���oڡ��*�5 �b��q��B�z'u�!������W�Z�vv����"�r�dn�(�M�s�(�_bt��to����7�7�L�Ct*[�a�����j�_�ٗ%zH����=P2f�v��7u"̠��`���ݫ��wYͻF`��h��o:�P�x��P���y��n��yʌeǵ�Ȉx^Z��L[W�:|��kѷ�6v�_�C�\�m�1��޵?:w����M�x�����y�"SË�@��=���/��Gm�,Y�����(ٓ	���UHW�6�%��&���r�[E���͞����8�RS��w��U٪eT�^�A.n\r����A&���K]b��ZQ&��y��<	\Q\���*=b���x�"��q�p����&�z�Ja��ts�v.)��s���R��ݲ�ꐸ�m/p�N1���5%!_����l�H�2h�6��Ƽ���4_H<ts��@zp�C5z���׭��+�����'6\���K��}j��Џ*�T��gmx�dI`��{��(����&��%�]�+�:�#_lq_�|Ǥ9n"y=���]0��Y>Kp~�q���9=�Wc	<%�n�b��<>Vo���B��״�ʩ'�Y�:��#IQs��|��JH��R��RS�3I�>d2�d�t��-�`�U����-�|���Բ׾��Qs���]����p��B�ų�
 P�2��M5��~{�Nz�<�Ґ�kc�Z΅Lͭ�����t���<��e�p��r�Q���'@-B�rsN�B�X�5�7k� �k$/�e:&s�3 �m,/�'ߺq�C�b؃8����}Q$�x��u�����"}��rĞ���q���*��e_||��!���c�:��ڢ-6�*R�7� �&�w�Mz	!H�޻�@BQ�B�H�I�����3>�3�7*�ܳ��k��}VҿB>�M�H���l��-�ݱ�Ǡ�Yy_���Mղ�w���HWQ|<S9َ�C��	�ɿ$^�+!���~�>�G���?G���Q��k�ҵ�b��$�ޟA��2��EmҘ:��~;n���?� :���[��e7ɮ,��u��RJX̷�&�7@`���p$ftr�(�{*B���X� lV1�V���/N�����<�U��mk����U������?ʔ�,�S'J�>`Y�V��q��n>(��o<*�iW��!�Q�Ǭbp��9�����4(�����W�C�ʪ��s�0c�j<U�������d�v��5�N�C*X�{�O���37�I�0S �I�$�t��&J�^��C��q`�2���!s9@{ǂ7��P3��z�|ː�P�o���4�𰽑6@^WNܮ4�ꊂ{A۳a�f��C<H�L��d��=]�R��0��4����]\o �O��T~����܏mϳ�3::8��O%q��x�M&��r>�%S֏L�Ǵ�Hu>���&���*Ȕ��E�����C�y`o�xh��^*�8�r2���F�8�a��|yVue+@UT,%�^DR?E�?U�U��[y�w �A����o��|��Eq�[�����-�F�$q�������I���lBZ���c�2�H���$�P��1ś�ψ��؉7h�+�6/���M��o�6�"?b�	8;��P���U����>��B�涖&����M҃�XQ���D�^�l��И��+��Y�4���3k�P�\3�g �:ܿnb��> �)���@����@o���>�K�����㾛��n^9��>�<�R��>�������G$f4�����6} fHž���ɗ��s��?#��K�� �釟)�}�h��q�)A���Rڳ����e*E.����b�ߝ��Y�IN����oE*Pr���1j�	�Nr-XF؏0�����˗�G�a>����+�N=p�/i��~3i�/�O$PE�2�. e�;Mء~��_LQ ���yW-U�VA(���ϵ�ԇ�u 8����J�鋁3��4�U!�F��=:ϥ�<E�\l����0+�b��ST��9B)�I	���So�I1�)�˖Y��)P�?p*�}~�Le7C�(@&�A��p���`���v:�`��Dڿ;�/��I�a{x��He�M?�|P0�[����v��hw���#e~&�?,rXrKd�繝O&�����������!]a)�������͵s[�~&~e��s#<E�JU�-35���G;l�Z���:R�N�g2��=�P}�-<U��?D�bI���(nk;���߳N�;K}f�
�=�Rd��웖*� ����
��Z��/ܚ�a��[�����t�Kb�
LѣB8hH��Te@��.�>�=��&=��c5Yo������[՚c~���&�L���s{u�b�v�n�ƍ��Ҽ�3&��U[�G��;p��G"7����^h�+h��cg���=u�:�!��+ �{G����0���_��E�ZqX���B��t��&�-����MY9���c$%�����ms|�-���pԮ9m�N�����O�ٞ��lu.`���]@��,�F+@oe�πs��^Q�2<�kl��\V0j@�D˽b�A�]�C�ē;(��.�� \៬^���#�Y Y�=�IY`I�0�8D��Q(�Wk(vy-��gcS��c��ǿ���	�n͖a@��Vx�4���_.��r{wa�G
�9Tg���Ӕ{;�]kg�Ⱦ�#Ok��]�?�H��/n_��z�)�A)M�e/Y�� �W_~� b�#E��Br���^���iC�ۋ�����K�*��#�5�e
Ũ�y;�+Z�>�;{�}
��\�ض|U沜��/A[��O7��:��ˍo"�?řIvx|\��8�sp���ӂw{r��h��y/k�F�u�-#+������?���]��`���l��(@���qk�-�/�f��>N3��C����P5��m��$��(d��&�_v_�6>�-Qx�#?Ӈ"� f��2?��@������R�O����-6��G�Ҏz<囒[S�Ml�P)-l�y﭅
�x���5���5����ӴE��`��P�3�fQ���tZ3)�{�?j�5��:=2�ۗ�����$���"���Qmɏ���Hqg�'xz�o�!���p{T������㹗�*i0�cR�����B~F�/b�j&B��
�1s�l6K%/���{/��.�˵���ޡ�Hma�cw=�䠹-�o�`�������[4���)6�r�v��U&G�����d�w��Ӷ=��L��������P�ǫ��^孖�����捪��B��!�!��)�3#e���$����)�����	�@���EE��l��U�����J��.��ɏY�5���H�xv$q��s���	G���/
z~u:�v8�N�6g_��O���:����S��|��.�3�G���ƿ�鉦,�P)Ga����v�75�b�0�.���/��T��?F�f������I�]L���pt��Tr�VRO�i���^���'9ps�Fzd���Vuv�`t���I �ǐ;`&�]�+�m�*<��ɝpL���)��1r��ք�9��T1�������w-^F1�:v5�}W� .�������Ԅ-Ǻ DK�w|-;�d��������L�w["���$XP����b��NT�l�u����f-W����<)waa�-�����r�����oG����͡�ѹ�8�Jc���O�Ʌ�>\3��WEpy#���u<�VV�Z֐+yu�L�d��\f[�5�����{7�(L�[eΧ�����) *f&Z4��c	����a� �Z��]��_5��+�m譸�eU��x��jU�mN��t�G6~x?��4�7ذ�-���\���gǦGK]�0J"b58�R�!�e��1��>qJ(�a��+��@n����Yd|����eH���"92��
��M�V��:;8�Gm)�W"}[Gv��Й�Wm�s���R�5��$��?4��4�ɧ��)�7�~��^R��q��^�Ԣ)�~��|KU��\gcz����6� z�����^w�kJ5M̈́��E�T~�$$h�\��M�Rs�2�T��t������b�C��KkP��W�3�r
r؞�Kn��[W���O5����Z@?��1���G�T��T4���Q�Wbrt�S'+<���TN�,�Ww̽�d�z
���{R{�[�ϙ�i=�1l���3(���:�t<*C��z�9�� ]됴B�4fYi��|�J�a�tL�l�nl���HU�����b*O,�:��m%�p���T���6e�iY�������!����*�g�}o~�Ǻg1ec=�'a��K�������f���f�0��+���)iL�.��)42�ɹ��K�o[50�-�Od�fa�:��!^Ƣ���>�Ÿ"8��$T�C;�d�0ʋp�7�|$�^�Ƣ��@V��v��$x�|:��ݼ�Zl�q���L�S�����c'��E�,���, ���Rk�{\b"v�2?^�-/��*��B�:Z�1���6=�R	�6[e_Y�-l5z1���%jNM����x�❪WM���.�Rף���������[Xƃts�Q �YfZ�G�����((D�x�{���[ g1�Ͻ�W�G^XtL-*����G޲�	��k�)�FBBM�`T� ���^�F�B��d2��D"���V�3������Xf��m���sRM�6�Qg(�~�|跢�����`��S�/+���_�g�qz�^�k�6�q��6f�9ڦ?���n�KF�E�����"�V3�M6Ƭ����5 ~@���Ƅ��Lݰ���{/ÜD�n�(����}R�+�<:�:+)���`q�&!A�����lQ��p��4�1���3�G�� ��$�)�#i�������?�^;�.�%�L���C=�Z�KĽz�`��W��������1����"�i&�/��=�;��r�(���Z�r�rD�'��x����ld���֠��0 ^�HJ��І>S!�g􆟇�����kˢ��ֹS.>��}mm5�Ts��q6�	ڪ��e���Y�������B�G�"�ٶ����-�9O�H��8�*;�'��S���c���'[g�^��I��Kޫ<C�]�UW�M׌�t)��p����0��б������ !�J����Mt|f�ӻ1s�r��#�zԜ̖���&�Xo���e�B]�<��21 '�S;Y���e���`�I�_�KV�1v�s8v���,9�0�Gg�[ ��T2���?{'����Ud���S�潭Fi�bI�]�����2KAb184�k���W��0�km	��2~�|��G�ZMl�����+Od��<�1�hj4��� ��C��C�%�!K��.~�1ֹ���5sȷ�>����Syk��i�c��Y�$���\�?�א�����p�&�%����~��㘼����G٧1Ƞ9�� ���<!�17�Ԏb�l����=tQN��5�A޷�?0�X?9ݖ,���|y�޲��P<$�Bsi�GˋG��O���	�����_�w�m<�i��kn���?�I.�:�G�s
�\r|� �"y���J%��C:�j�a���6 qϾ����bk�t�蓲Wt��v�-�ܹ1Q� f6s���8gѰ�@�\�����!�j(�Ԙ�o�쯫k`F�4	p�Z5u2�@��)��c>i>M�q\�薦t@'Ǒ��*��Ӡq�����Ds�1��?)M�>�Ǿ�S�~�u�T�����I��#���T�R4��Nmk뭸���2@�qs��xo����uGM�vY�&�&Ɂ��Aۧf�VР,���D�"��tb��gz*r�QȘ���/;�t�=�^���Y*��/-;Tu�@w~���Z��o�"��j�{��.q�T������Hj�sm���):��y��I�:'q;xQ�gx�6�KBB����j�I@c�AK"q�qmY͸�`)q��w���m���Z��+���E�)����+��l�����D/�����D���{����5;㡜��=j��L��s`x��X����V=-�G�K:��עP��\>��D��o{O�ͥ
�B�sF��uD�������u\��J��j�y4�q����`�!Y�t� ��X`(o@!턄��6�̈ć�9��^\�2�9�;9�JFdަA�W#�$��9��<%�.'QtϘh苞4�����J������vtp��ZZiO����J��D)+Gu��g�>CY�:�apPEm��cW+��*�r�w��ov�MRg�����g��l�]{G���-?,B|Z�}�xWRXj?��d���Z1�7�Z}�f���dΦ��5�� L~+9o�|�*h�:���ţ��F�;E����q���@�Z����ՋШ(���)z����'���X�`��T*F��Q����k������N8/�兼@�S�5�Rs�bL-�����|_�Y���5�	@�j�'���p�'�x̤��'��*й�Ҳ���z�\޾���� �k��d^�c<��jQ+e���Gi����F ���h�|������Xc���n��
N�v���_A�Jʊ��b��z���TY*�!U����o�7�
���,i°{���s��r�7�<�}����σ��Fy}��,޺��P��_'"<�7%�B��d2�:�f�w�Ռ���o���z_���oؕ�\z>+@���C�������ĩ��n�˾λM�+���u�;�C�\�r�'�ҵϰw0�����t4|�Nv�MU�g��o�^La��!yE���$�dJ����3���Q������Ù!W��ufF�W�7bkYd�M��/�?HcȀ�C#����a
.�vc�TS����.�u<A�$E�K�|[�a����t�N�x��D�$�ׯ�m#�r���uV���f�L�Ͻ�Ë4�[� ���Z��fa�s��y���Y�9����R�����c��F��Tc�|Q3כ�vʏP�W��<���JZ�xU^�n� �CC��T��\��v�ja�X������(�\>��C�?U��B�Ϡ�2�ɬq1���8��%�O4�]�B�M���L���TS������8�j#'��G�
K��@@|Hb}=X�"r�<��x����Y��(���B�׎��h����0�����>����P[����:ɹ`�٥�uV�f�S�3���K5�N�������\���[Й�����s�dϟ����{Y�97�C�e8ESQjEz��GC<���Ի1��Q2:�^�j`�����җB�DBJ���9C ������Y��;BB5���H[������Rc�.ǳp۹���튗��I*�����m�/�� �$�$�_�~f�5=3b\�$�!@j�t\��e�}X�<>j���/-hTR��Zk9�3�_k�<¡P�*�A�����W��឵,ܥ��m���	�<g��/l��=v�����&��ǧ�Y2��F#N����cc���z��e�Aj����w�^�1����������H�E~���J��Qfe�c�z'�_
�6n�m�t*�ϕ�"?��7_H��'[��&� 1�1BV+�E��X*�3�1�{�wPg
P�3�ظ����Y��wj�L3���.)k^ 8ܐ��'�d��0)����W�X���~�B=UH�w!`�m�Л��2�����u�E=͏��`���w�?\�!&"���R���=�aX�p`j^����/��=y�i1#�������R�îw�|n��JY��H���B�������;*�%I{��._�F45�H� 3KgB@M<��1������o�,k�F,�'����^ל��uupe�c����z��tE��_W�G�^9*sv]ŗ>��j��ih[%ǈ�AM�?|ȉƟ��/"/�obt�^�G���$� I���k������l���1.� H��~5,@>��\EOl�8hkvђ��Q������rW�����6�~�����"{HU��Ա�_Ǽl��/~�YP|�y�a�.���r�\�8�&7���F��C�b��L�c��B��?Lϼ55u}�7�T������}N�on�w4��U���r5Y��ӕ��y�C��G�]��i��R6�{Rǫ���	 $3�	�>EbF��vc��=I� FYXȞ$jg>">�&�/,ɓ�dz�'�t�6����X!�'�ɁО�c��u�!�۬ ��3Gsʍ'���Igz�ͻ�o�ϟ�7�҅����_�a��ˋ�rp�*������������Az���z��\��W����"�7�w}�]{��]�o�1Zd��ݾw0ފ����Kd��G���a��O�����;E���+y�4�OAE�jW"v��Հ��Ý,P���(�^'�ߙw���/n�x����uե�����TVj{��hW��=#W�J�]�t�H��8jȔ�38��h:W��-%�s�>���w
�k4��M��u�#E#'�Υ��\��p�Y�w��)׼�+>~L��5�|s��{_O��~�����ޔ�`��tv�1�a��"�}dܼܽ�u��<Wީ��D��yw�Q�m�U�H��0I��)�}
̔����$��)����?����V����a�Z��ρ��ЁZ��o��9J�8���P#�=�+e�?�-,���ʼ¿���V��5�8��2����7jtO�u��9w��=�Dw��)K��r��C��|�xX�9dِ<BK�|h���E��S��6��	OW��ٕ�~�,&T>Ǆ���)�nT1h?y��~j<�E�����(84�����'�\{����\z�w=D!���}�S�y��q��9S��:�s:~~�\ܦ�<<����ᗵ��,��qx�K�~��)�mS���ZۤmJ�å��'��7�XZbz�&J�sBH�W�(q�q��:��v�<�{\�qN̯�Ӡg�/�&n��|}�BM�\8
�!���_��i�|���z�V�Lr1ն�U
�@+��|�襻�R�J�UZ8�H~�(+�ԫ����Mq����˝O^�ɝ#�
��<K�C�F�N�R֎�z��͇��[�}-(�X�2�G��8k;�`x�-�X�4�a����"z:��F:覎u�n������x8E�d�r~G��__IB�|��M��¾���}J�#fn
x��hh�*l{��UƑ/,�V2ޞT|�י7���N��.�U�	��K���'+[��SC�kä5��s�H6�99����E�[�#kq�ǀ�ʻ�}�%���+&���/0�`�T���K����g2/�-zuaf�G�p�ɝI�~�D6�&ҧn��=�Dou[%d8�b����A'-Y�����i��O'FF&���1�G�qi��MY>K%ۘ��eb�43�����G;�Դ�) 
��T�Ձ���{f�L�^S3�1�����^ٳ����E]�@v�o�l�����L;U������N�uY�3o�_^��<\��ș�?����-�#a�lB��/����Z;�����-��o!�6Э�����|��G���U�Re��6��Cy��=��~�=����x�.�K=�����7��{ Y��o�`�^`�-s�'��+�h�V�w#s�O����&�t`�]���S%��b&�Y�Hf\*�~��x?L�u���CV��V�ʿ��$�
�|���E�ơ{��^JX�i�����/��j�3�a	�����|Whnƭ��7�^��~�\��l�Ա}:������R��G�yv��sg���\+�⒚�2�{��8�{�5�U1ҵT����Q�g�*�܎���0hϺf��0'�v�j4_f3��߉<#�k��.3Y|x�"<�a^	MS���!�%�!���A���&Ψ ��<ǝ���\<B<3�u&.��5�z}�hUT,�b�[{�����Փ�z	��ƶkt�^�L��R�r�s"`����a����������VkcE�U�ɞT�4��F�4�(�-7��P��ʛɋ��#�����M�N'F�9�b=E����iV���O�'�Whd���Rd|��_��o�?{���z�;O���/_��ys���D�	�c��syq�������	��W�Z�S�����r70��N0�㡉���7.���{ոq.#��Pnaa�o,��O�.�kY�Ǜ�A��;��FF��������K>�?�f���niK�U�0��z��M���'(��!D|�!�rr����;�Sv���5����G/p���)�]�#�טa�O�U�/��{�u�z�A|�T��W�i��_�up_�����I/5܆m,�/��&B�y�)���ng�g
hP=T<�A����tU�ӵZ���R��Uap�Wk0�_�e�prm�!�OQ�(b����D�!���̼���NC���ON�]��w��N��H�� �6Xp�W��%1Q������Gk���k�f쭪Z��}���'���朷�#�Ѩ_�Y�5h��;���c&5��å�j�s/�#z~E���r�}�R���إ��L|���R`�_LJ񅓯�4�1�Mΐj��yt�}����'�����u�qH�@f(�2X��x\�� ÇAnhɾr�&\����@9�?��'�2AwG�u�=i�6/���}^b��v(w�p����)#aCX�K��/��lH�A�z��w�~~.��*�se��a��Ov��%��Y��%��\��yO�;?4�t��F\�;#HH�$܇K�G��l�57��5��Dq�[��]�R\|	\ܹᗡ��R�+UXXh.\P����jt�h"mm�X��O�#��R���Y���Yಷ�4�V�N��7��y����
�HLQ��kÔ�s����<sΩ�]k���@O��t�L|@f^|u��{*�@�|����Û�K"��3I;Z��tnd�]iG�HK�~"vX����Yof�V�`��>ãmö�z�o6�3ԛ���|���kl�m���j (8�Dr���-O�9�\�ş����+�}���"������%4*��w�j·�,�jځdu�ų��ś��A��Ė=�3)eͣ�g�@�ҙ�Q�����*nf7�yi"� �	��	=)�F��c2=��T���.a��ͺ{�֬7���z}��������d
:���N9�kM���y�T!9G�a�v�Z"���l�����s��sV��b�[��e�T����7J�	o"R�Q��q�Ғ�l�L����l���p��9�m��cQW�خE�d�C�ʥXe,�&�����1�[�] ��c�ť���1�.������9�G�5��r��<�S���5Bob��\�������G�*h�ؽ���$E�4|g4�|�_���O����W��ZɎ��v5��I����K�5�nM�,.ܤOXV�-�"M�:��K��^im]���oLk6�OѺ&њ�E^]���v
<�����Q�0���8΢���r_�qy�uP�H�E��a�jQ�M�|�ae����Z�ꚠU�<*�}��P�ꓷ���c�p\6�3��$�T�]��1�
&ϵT�������-���y<��-ɞ���<hC���=��l�}8Ԟ������Ps^@����[�E�a�C�c�)�E����+Q*fhQKI鍔�����R�����7`Xˮ����s�	�%�&���W,?���d	��׹}.�y;�|�ʕ�#6����>2�&.���.]�,v����R984ռ3��Ll�U���^h[ZR�8QgӼW���P��`�aJ܄ Ԝw�>Y\�u�D�K�Jj�<X�6s�(E���1�Q�3?;�$�\~��yO��d�C/F��ؾڧ������R\\|�H���{���ĕ����ə���j��V���p��y��]���skf�P�߄�7�x#tu|¾�J���t޼ɕt������}��v���S��r�S.P,�<p�^nۡ��#"ϔ��-Ҿ�5�q���~��+i��+�y=�5��N�K���.~�|��q���dԣ��W5�\zFjM&}��#�[�Ϝ�>�_�s��A��-�����S�(��d3��!��������	Z���K�$[���z87i�:R{(/�&#u����nPL�u��]<�5l��]D�!�U��;��| �v�M��"Gz���u�lY���"�k,P�Γ�e�����\�K�"b$Eu��Ѓ���>�e�xlB�e���z~���ĆϱY��7�:%z�Q�5�5����0�G��Z��H�W��%닪[;��oY[���b� �r��x:�DM��{K��~��tw����-���v7_}�8Q��Z�u	��� )�S�%i�'����3���n�\�~O����(�1�!�[1���"�p=f =��g)�#�8;{�*Ҡ%b]dѽ�K�&��� 4K�oӅ�o�3�<��ڐ�	ҔJt��c��bi	x���0��i�c�QM@E�Zu��hq��ȣ�-����QN�쯳����'g��{{�Б@�bݴ4R}ass�13��X"�G#����=zNC���-X��.{��޼��J0����E����ľ�x]������������.�=}��YX;�u X�����"�U����r��{��jr{�y@��}��"�M����`�*Ҩd\dz�1�V;}�#���mk��P�"Q�B.z�N_��b��,�z�|�u���{��ɣ��\�`/���:i�1c�D���}d���:��Hޑ�?��)��&m�C����
��%�a�ez�cQ�N=PU���W������I ���8}��.���kbRv)�I�:�J-J߼�x��ƙV���~O��w��^�h����ar����[��]���3��\��-��"o���|t6�K�)+��SNy�;NV�FOX���kdW�^a��嘝��8��h���x֛������4r5�G4{{���0.K}�y0
���Dv:��)��6aE���{^.����O(���7zZ���a�Z�h�̗�w�n=K/ȣ�*);�>������Lh�lx`�6�4<j�f�}��^Ł�{"�Y�����S���)>�V�|�2�Ng-���~�?-�1�j	_}5���z�RC
H-R�����3�H�!������\���5�I�ram�$T.$̻ە�	��=�k����2<"��(�`@����<����s��1��"�fQ�<�=P�;���E��+��>s�����q��Y˙�J�+�,`S�fF���>�z)�o���]M�sa������]�:��v$�W�y���̑���;�e�+WF�-����Aq[[���د��`&��>��Ɂ��r+�fҩ�t �ax�qݨ���ˣ$X
�۹�~��[�.5���nk]�e\�.&���.��ԃ쟞#�����gpš㵦�]�^9��4E�����vv�
��%���(/c��d8'֯o�$B��r�M���o�5����܇��� ��	�2��g�:E\	x�^� ���S��;���ۛR�C�t��o�U&��ڥ�:�y��l��mH���Y��|�_�@��w��g ��PU<�R�!D ���Fh���S�醊2DP���]-A�<�~��T�����d�i5P�b�#�:������\P�u�i:�����T�`��J��{6��Q��/��B,,ު�%�y�2ղNrjN�J���f�����G�wD�Q��pA���4So�`pP�J�8M��U���)��x�)x�1�*ٳR�^��pbW�B;@h]M�~�RӇV�\VnGݩj�7������T�fB���FK%����<m૵�@{<23/�:�����9wpȚn��$g=�d<�)Y��PȖ\�&輇��G�I�\�[���Iz1����u�~O��Ga���_u��\V���#���yT�a��^C��Go���ܘZ||2R����t5�;Ӌ!j}���Iɩu7��j$Δ�����h����ڛ����Pvs�������Ռ���Od��l�h\hx�n�%]�yT�4���f����K
L��.L����J#�{e�5F�2�c� ���x�Q �@;߯��9�6���s����9�܉�Ȍ�9���ɓ	�HA��1.�yKI�*C���4�"m6���(@�Α�ƾ~���[�4��ǫU)��86A��K��q���!�ޓU��L/8�2�f�.��ʮ\�b���fȣ�F�ߦa6Y@°���)d|܌�ٺ��ټ���ȵ��qz \�Ih�|�u��1kve��-�8D��W�M���ApH���j �B#1Aw�mU��:�����lSa �e$�1a測J����{���uK�,5oD\�(�NGR��/���c�Ć���Yb�}��4vG�V_�j)�4�ap�U�6(��(����E��|��z~�ީ�����]֧�Ԩ��T�S�ĮlSĔQEg�Q��
��K���*Q<��_��6�>�w�º��V��#�L��������~U�]4M�ʹ������fc"r�_O�ݢ����c������@�������&'��Y����n�N4�h��G6�_c��Q�1K<�ѣ�v��)Ϟ o�E|ջȈ��DB<"������}�Ѹ�����V;TF落3��n�\����V����|Y��Xʨ�[�mZ�0�N1��C���/RԮ���$��mw����o�,�`�� H�l�J�:�XtV�2R�͔���͢fiIՐ0�$��޻w3�N
~X�E	y �^>'�L�����ּY��Z�2u!�g#{ �|W~��y��N?֤%5*ntZ��I�=�{�J,�����/�Yg���Z������Y�󲃆��0��ZT�3��a��(T�Ns�7 �·}s�o�`�純Í��O�����=nlėEX1���m����j˳��" w44�p�����y�f���#x�B[�_q�H���ȉʗ�yϻ��¿QLv���'�@�E���� �x��P�$�/.������8=�C������n�!{' 3)�e���$^�lC3|� om|�gNę5yN��ȑ�G}�G���+^�_:�xQܺ��r������w��Sn��
�®v�_x|�S#�O[�� m!�~l�#��
;z�: �+�����2m
(|�
E���'>�@Ƴ��� B����n��V���7����[��
>�� uu�	Ⱦ��w��Ś3Q��6Н�Ǐ��k�[p�����!{�P)l��n�=U�Q�'�����6�5���1	����D�\حpFFd��N�D�p{�����YA�s�]tr�-�m狁�(<֬��Yp'"Y�k��E����t�K7��h�m��DSsu`���QrA�� !qb��7e���K^cb�
c�ס��f��8���䚨����y�XO�k�D�^c&�$���9g���F��ό�+���J���%���kU
��+Z��G\NzU
�TׯS�pGW{�xyƮ�ﶉe=8X[�N������c����[�ko2�ʔ+6�/�����ơ��A����������Ts���j]AY��P�����M�����V���BX��{�?Υ4-Ш�F8�T��-X�f���ə�W��T<�gZ�u�w,����o��4����R��$L�q��z��U-��W<��!Z�0d����O���JE�B��	��룙r.�����fb����'< R��5��z ��VK�%x���I�ȴ�C�B9@{��؉Ab)Mѥ<Y�a�n�L4�O��ez�̉"�,��&�R�.�[᝝\=L��?UW�)� O��{ ���
�b�r�\��8=�X�B�wm���*�>�G5�8�\�F�B�e�J��	���W�Zo���M���
�J���hn��-n7�����@e]�t��K2�:�s�|�a�3�߀a4����UY�7�]@̯�Ǔ���e���'@�r����e8��]� ?���a���-��YF�Ts���l�t���seSU�D�)���]D�O��Z����;��Y�;S&��.����P.n�g9df���B��A�]>�%Q�!�.��:~�ĭ$"���$��5��ȿ�����6��=4@�[�J{�c0��1���&�֢�!N��t����Y�2��}^��D��Sd���c��m���I����	��m���T������_�X���s�Q31Y.!�E ���^�6/�n*ve�]�W���::e�1�'B��/Rj>ɑ{Pq�aDR���`�r*������a¤e�� �
Z�C�ܹhȳ4�'rh����cdT��%��� 	��vŰdQǒ%^zn�:���۷�k�P�Bñ��DZ�a�zy�Jqy����̀\:x��|qh�Q�a-~B^pqQ���U�*D��ZB�����]�<A<�u,�|�pE�?^�q+��W|���qD��7ؓ���1�����X����U��~��^(����-�5LSĘ���A��̲�_\"��b�)6,J��^�����m������S�O9`!���gY[�zf��,&˩����+S�ri���wv�h��q%�~�T9Qz�ʕ�]�g��V�7i�um7T�&��R�~���������/h�F�܀���΢ �o�`©��G� ��3c�3��^�S���D­Qp���&�/��x�e��&"f��u	=^Xx@�P��x��-ډ��/�.�������Ve�����d�
^��:�����"��Qin����/G
�X�1��"�	���&)��زo��o�c:F���yq��߿O=�_�c���vC'|.�l��5�.�ދ������xmYD�[��󘘹 �*��K�L�jγy��_�����#q�*����}?�:��g�e�p�$v�A���!^��6��4��Oz"���d�Ix����6��'q���5Va��U�E��Z���\�m�4b��&��˲�&����Ӳ[��z���R�6��1�$3�O>�J \F.75?x��)�ۭR!�D��9bΆ��G@k��G��������˜ �~�⪎;O}}U#�FuX�S��w��kI�26�H��~".�X����ѥ�.�1�/hE�B��
��?O��xd�Z��X�Q%�������!۶m_��n l���f{zĆ���ę/�0 h�xM�.�*���/��c��$j��2�Dap�k�Y�T��J��~=�Dn��d�E�R��b��o�.zC۲Uk,'�J�*�o)\qH%v��C�(����b]s�.��M �p}�+��~��§�=��ɋUV�@�qL6�Y\ Pʌ_�"�CfV�@�k]����]�r'n����~�=�]QVAR�޽��;���	|��������rZؠ���"b��\��݊��5Pm�::��e�p���!�r�+o�����L��m�{#�(�5�A��~��K_�0���AY��,��F *���=��<�0 ��{=��ň<�x�c�W�5k��?�M:K�(�Bg�8@��F$�gέy;z� �	�M_�Lk :�����ΕkRLP@rg@e�rF�	��?T�[�(l���Oqp�@>�M3+�iC����%%�=�o�,�ۖڠ��uӭ���1_��8GiZb~���E�q>U�q�Xݑ�y�ö���ӡ#�f��U�o��AgW���Q�A��9ݰ�ػ��ؑ8�R��+�=�'Z!R�d����!�n����
 1J���F���p��}��<���mD���hf�����_��
(��GO�]�ӿ'-��<l��#�~�VR�p�	���0��N��s�ѠjT+��f�j|���[�<�g�Z�T"b��d��o3�`Kl0��P�Ȉ��q�;�:�p��5t��X�
�������D�lU�m�ʕ��L�咁3��^kŀV�_H�%�����ߗ��=��
�W5��ԧ:T4�#�Rk��|��)���I�z��W�F�e/Eea�;����Ɉ
5���Abު~S�� �![������U`4��a4�~��a��á���aZx*K=��Y��"{�}(�2�}/�E(D���}3B��o���e0��0�{��������Q�!�����:��s�78���XO�� o�k��&�m�L�&%�bx��E@
LO�2��S�>��e��*�`*N�p,g�*���X�	����NWY�|m3x��K�8�:k�Y�2k�W>c��K����Yn.���r�e����_]\- 8g�lZ�l�rY��f��DP�ŗ<�T�!�7�j@��S��?+p��E��4�}�<��c�&��C;�Oޚ�L�w�u�����Ty�d�a<�B�mAD��z���bO��{�dW���75�fDOE��Z�,��S�>*r[R>��G�I�̟-��;6�j�,D��Ƈ�?�kUA���/5N܈ɛI�CyF�4i���W@x������rv�N�DT���S�v��u�?#�?K���˿y��\�c�/�0�mO�{��Ŭ2GhmO؅�xTp��*I�ꪫ�J'�߿-J�x`l�
�y���CR��xT�_���H��2ۑ��w�=]d��VW����5�Ɨp0����������D�.}��:~�;cj�D�jA����!2�4�;z�ZW0�./�����&ݱ,�(��N'
&�Ty�нfr/ h���P�\��u�$���ð�������l ,�k���6rŤ�M�:�A�h���V�&}S2
�Oň�L�~�67�ܙ��&{���&.�k@��A&Z
e�\;W�g��}�M�}�*�O�z�4��'ގ�Y�;�e{O-�x��<�Fl+�;�\�l��q���M֜���rl{q��>��<Ϊ�lm���^���T��x��Z[���сfǇ(�;딡��Q��<����~a����S�녪�_�o���v���QS�>;�c}f �N�_��(<�wQ��2���4��S��gO���4�|6�N�jffS���Ӗ�� j��P������O���H(�aiDۻ^{��'�v)�rax��� ��g;�@<����ɤ�-�ų1��:���D��gӍNdp�2��FP��y����~����{-��t������Ys�
M?Pb�
4%��+Fi���� ������u��S��ޑVD{c<v����RHQe�N~��]�`�Fhh	 �4����W�����"'g�G�T: )M��� ��۞.k\@��z�����˕!G9Xz:��-�����`��P2��8������uۿ3}�;��C/V�;Q0l6�
%m_����4�����i��y�l�_��MY@�O��L%U(jk��f��ƪDH� �E&w���k�τ��y�$	��/e��!��$�;`���ߌi�}h7��bk��2d'�����Degd�M	=u�����~`|l��k��%MsI�:2��^��R���b�]�>��@�{ÿ���*&nyHc�1<�;f�����3�w�p&
G��<��gަ�ol\�#��'o~�[��B����p>�]�WL�觷eU-*��{��V-��8�7q���HĖZ�o�oZ5�1��"��b��·1$� G7����b�S�b��~k=&�fgh����튏�� ��}]*����ae���C��fӸ� ؝ǆG���Uhpp'�udqh���|*��EH2�Jum���n��H+�v�	qf�G^N�]�n�c#�\-�=�/�e���J�x�Ke�t��ŋ�=8['��{����1AP���R���P�F({�\�$ef�B��j�*�֩����n�$>ȟ�y�^��A�����qk:�������N9�7������-AB�]�����o+�mY\�12+s���RGJh��a"{�_�"�5�t�_k|��mQ��м�������"�P���j�>�L��'/_�Q�5�v�����L��t�}�E����`q������p�~�#�T�K0�s�P6�]?i���_�[g�e�m�	|ۍw!ݧD�a0�j��3tc�������+�Ҷ�3RXq��@i?K�����B�;�Kp@ArcżMZ�ٵM5�Li�l״:�M���OI�^M
ˤ�%/�]�6�;���c����h�����U=��k|��|o��Bت �8Y�Q�ȝ�9w9��Ot?�������f���L��=���2���u��WP�C�fs��S�t�	+���4)�A�ȟ=���N���? ��ޯ�đ�|S;XAp`E薝�^��h�����6��6d|z����"��sh�'	�C`<�Ic�z��[���:�J�7�����e�@.���fגʡ'Ul��~n�m�a�T���!��8s����5÷ww�Cl.L���3�~�̍�֝���"����Ɠ)�M��ĝ�}4�g1�ΟB������k+s/l�����,U4+��Г
(;����go\,dC}��JkfϽ�2��x�c0��u�Z!����}��לۑ�q��N�}$�@n��9q��&��f0Wkg4�&�d� Hjʞ̱ޭ�g�:�U���#x�R�b�@R�_�boL;E=3�}_���q��z������a$�k�����;�J�]$h�,�}��/,s������,¡h}��im��h�Q�E��##uzXD�SV�C<� �����{�K�
�B��G�v���pTp�~(vA�~'����V:���� �H�-[�
���K$\RD4]G3��i)���I*�9v^����V&l;eӨ\�P�N���,���W�����̱��w3�ȇ&>�D��Tj�{�_��es���8ʽrLɨ�@����5�7fN����ߧ�Z�c���.���{�YwřW�D�_��z"?x�o|��:k����T�{1�1quU����
�t�t�Ůkw�ô\�2 %�����"G�D(Y|f��\�-x	����L�7�Y#�����nH�}�����7�u�NO�?ɦ���n.�n�GX��|��?�+|CH�.�帕8n5o��#��xaҤ0���h�Z,`NG��6i �~K��ȱk���,���Wp$��[;�if�;�'�㻵y��ˋ��T9�O�n��Uy�\�/I�q�7�7#��~x'-q_� �������� mP��z̀tO�P�a=@�+m��%Q/;E�仚�uG�%)q*a�+�����|�WگAu���V�52�~~,J(����m��Z�8��y�Z��w�%�DD�����`���bP��ڏ^�#��LXS�bC*��(S}�{��Z��-�aPЭ�{<5HV�<���?��YE�l�ՠ�߰������q����p'+�~3��&�u�`��w�y�?�:��M�9��"���g�:�r��2i.���qB��(/kq	>
Zm?G��>S\ e��#ݗ��Q4�����P�H
&/�}W�ﱾm�g�F�}X��� x�+Ic�Ј� q �y�J����M���Џ��1A�C���'�f���@�i�5�{U�I�谥�K�>h��#%��7VP�_���4KͰ�^{�Dܘk�gꬫ��4#��5�/I|-~�pLkn�K�������u;Pt�>�p=q�^Xj���	叙���|���fr}�4X*�w�x/3f��=[�q��ȷ��
��#H�7���������b�[�O�ǩ�/e,�MC�Ǳ2���\�c�ᔂ�����U0 �"��۷�mc�pd�ww��x�O�CΔ9�y�#���⩍1s��B��U��n`ڕ'm��G�����;�ܮ��
3����4������vW�s�Q0�0?}Y�9t~Z� ��
^�	��Zi�PU!��0;�e >������I�s�E���4[���z˟��C��=Ȇ4�|;��t���V���� �=}��X�3"9��X���)x�@�B��'��T��\�e�^w6mfȰI�ӠfJ���ɺ��?@"D��Ġ�����c""FֻC}l;B�7�� �S￀��(�U|��oc(I���1���j���b���-%oqN����sCby���war TJs�f���}�E�wG�wu-��+`�u#6	�p=� SU�.u��Ӱ[�d��=��<GF��矚�8>̿'�Ř~�3����5ϖ_C`33�3�*���b)�c���;��U�ܮ�b@60ݽ�wD,�T̎�nE7r�:����v�v�Дs�ݪ�R}Z3��9Ȇ����t3���E#���&UA�R�F �(z|�7"�$��C#�C��0;?�	K����uo0~�jvwp��$4~ob��u����q_�p#�.7o~9�V�9�8������O2샚Z94�Ld��x�m�L*�C[��.b1㍂P�i���5?SO~����x��u~������D��^a ��}�*zЬ�j$�Tu���C¤��4E����̃���6�-dF7.��p�;�]��0�;uH�xT�	?��Q�j!�EF`��!�5B����aoy�y�5��%o����llk��
���GJ��{�p��lLk�����y���yk�P�JL�CI�2u3��4�k3<���}�({:nn�?��s�+�����v��Ĉ�/9EE:��9�i�ن
wCj�ω�L�t��?��^OHw�z��7��QA�N_�!���k�Ǵ�@���
�24��c�á:�@�$�
����VЀ�3�J�V��\�ez>�gyk�ʊ��h3WT�
�Nb���۲-��
 ��#��tԝ�!�H˫$�U婲���IO4X��Cx��_���jj�@7�
���C���� �.� u1��+��I?ː�;5�,d2��w^���?��P���d��ٽ��L�?��;U�I��Z��5TB�a�Um*�LgU@W��.H�cr�M|��K��"��d���ʸ�^�8۔�l�0Ɗ�'wH��pEuyt�cQ�̙㇯VQ��j:p0UG���3[c�Rd�������H|�ډ��v�g�݇�'��3����!�TE��Hl�������(y�߳��}�� �a<R��ν��&E�!�&>�s���iC�����T�c?ji8��x�S��ϔp��-a�[0�#⯥�&�t�H|�KM�����w%�l��E[!2~�bj χ^��_�x!͐q9�Dߓ�B-�ŋ����r��Պ����^=��\����A�CJ��FW��Ə�P�~�������/V����K,�
0"��]�:/ӻoG]5���Jy=��9y�~�\�v
���)����%dc1@t@��=Z��������oC᫫�z�3Cp���6h"Β���=#�Ʀ���P�;]=±�1y���ݹ͍f�,�n��akF�juP�~n�;���{��T||�"�>�:��:��V�H9�s��גf�oJ�|�޻��^��8���D{u浉���zu!��f��9��r>O��\��fǪ��cSq��V ���*�o1�nN��;@# �v�y�!U��1ШÖE�G���L�9���O|=T,V��(��"Cu���{M�ki��o��I�ܓ�H�ij��K
R��_���U1ij�Zy�N=�7��X:�}��u���C�&��P��ZbMC�a���v�f�{�|������@w���)��$3�������G�P�;rȏ��l��;�����]됤$n��r4XH��p�3 �ENh�S�����5V�N9+!^��u3�=wb���+��3��l$m� �/����f����Mq�M�"T�O�Z+�/�?�T�<d�i���ᤜ��Լ��S �V���lBJ�#�s��"�W�h�,ƹo3Ɔg��/�*�=�$O3��wmV�ZQ��rdo5S��31�����P�H]�n�fE��Ԙ:Pzz!���[�=b+M��+G�c>�
���L���1v+5߽��R�����I�Y���7 ��2Y�g��RU0vw��q�{@�4����IO� %u���90�������k
�9����_��D65X�b=W��~`"z����
�J�-��;wF�D��U<$Wޫ������?~-�r��9�0~,[T��I�>�B����~��ØLy<�v.O��3� м�``�$i?��(�����9a"k$Ƣ��;��/�%���(�2k<�g�!ݽ����$��k8��!.ZI���t_ۼw���Os�]j�爖��ȗ-`K��#��@��83).}lM:ġB ���&���P����+g��jJ_n��y�[�{���XZ�l
vJ���*�^.y���޹�[����}x]FJ
CT��rb�zu�q�tl��X�4����axȯ2�N�{�������2�E~��Q�)��p��e}̼��q`��e��ߚ�AM\)W�՗�%o��B���ڮ�>�E�Q�5��*�&"lt���*����=�����bD�5��襗^!c��a���M�2&�i]�#2��P���}޽�3�8�/�z������P���&Eh�F`h�{��z�;���aQ��v|����͋�t�B�j�����g�*
��5�h͡6w����{�ldRi���Z8����R��C��ۙ���������y��q�U��=�D�[�kg����/��C�M��D���F�@��m�X��T��`I訉�P7�I&��z�ҩNz����4B9M`�s�4r��Ft�w��Q���{w�3M���p���]ٝth�v?���M�#�O}���I����|���B�R��o�<�M�w:y^!��f���`��m�ob������M���(�׿���ļ�.0�sS�l `V���N��R�|tm�v�����xGSh�pA�J�@+
�Bj*b^g퇦�:��T���ψ�;$5ؾ47H4�*�����wm]��X�kl�w�U��{�7�����Yn�E��a�!ԇ�e�З3YM���^��s��-ڶ(θԷ|�,D&gd�K(@�����g$13�-�H˛dQ�>���vm]D�x{�����JV$���/�Nf�!G�:e�FC���p('���W�C'5�Ę��m���+�!Ƚ^=�sa�f���N��a�JSG��80H�QN�.iK���^16=�i�^�F^lye�K��8��Q�n�W�d_W8}���Ő��X��-K�x·'p�^a���0�>�W^om/��k^�����(�������m,��T�LޣG�:+�]��B��v���x.��h�R+8p�E�74c�<�(B��p����&N���F�D�4iH�<���?�q�=^⣝���L��I[qo��<��ՋW�j���j�%�0�d���[u)%S��;�M�l��V���FUA�_�W�!EJ�1Hw̓������K�`ZKӒ��~G~��1R��K�A�X��I[���\V�A�!���Mii�I�K,#�"�����{�!�̒z�o�9�*Z<������.��)sx u5d/�u׹�i���R��yk�9�!���bK>t���>���i 0d>z{���7Lv��W� ;@+�fEpS�tuM�a���
V�o{�|���s.����y�ʅ���w��y@��m|N8�h�~#6�Kj��uA��F�}O��se�)�[������qAu��ZumU;K�'�^����i��fU�a�����W�8�����sf���!	����������>D���46��};�R�rNfK��= R�$"�"( >kw��g؋���^���2-k�Z���ʵ�x�G?vq?X��9�∼aL�r��J���Z�W/��s�Q�	kSy�V��H���ؔ6��4[�?�U��l�۫��a������Tb��x�\/;Jٽѫ�zd�7�p��A�|�E��,���[�V
�W/\(X&�v:�}�,�/j�X�x�r|�X�E~�:r�Io^���[�e�:�^����NU�=��>Z��B<2:�tѝ�M�KL�y���E{V��J�u��HJn�������Eہ�ir}z�7�h�t�q�_�[�VY)ۛ�#Y&Lk�i�D��������U5��;�����4�Ë����Ȩ���]W��e������y�x��njU��N��b�{KD%�Bʌ�u�u>y�����r,�2�;�����t���й��}�������dM�k�zJ��A/����
��ऻ�+�f'�� �(�P�]���`������{}��?�[�|�<H#"���^'?n/I}�����Z2%d*�'oov�{!�v�D���FT�w澳I�����E��@�����ctI����S�y�Fs�&b�>��b������Ԓ���h�h�|�)�B���&���q�=���S���hT5����Oy�&>��ph3w��;�8e�������~c+��B]��������%��s��X�Gk_ȓh&����Q���b���-�<�H�7�ٰ�*�^]0�k��VXp/�XF�p%Q��:�A� 
-��bd������_7��[��F?/��# �856�i�i��R��񣯖���3�?��(�M��~0��טT��9�'���s-���+��q���$��>�qSo@m��yh�Zͤ�����NXӣ���Ub;\R3��|��߮�L��<�踼��U#yO/����U�1�/��	;���Օ��o;�*ήL�h�Ĩ,�$���5B�|*M2�Ɵq�e�pq�RK�L��!=`g�~� �Rp
�z�JP��siJ|h�P�yV7����p.5���N�>�L������h�F�؈K�
��c1����a7 �ow�Ư<s�z�ho�U���z�Ӡ�>6����v�Cm)y�,ŝ2���q�!�G��/l�����;�%��j�|W�d]��Pߙ{�=ڱ �ypu�蹮�k��^9�ZP �h��#�x3O�����AJ��'��m�$�7F���.�����4�7�t�/e��ʽ{F���� ��$k���;M��=No�G�]����i}`�[�I\����{(��qvS`*�
y��Lj��fq�vN��|�����K�m���n������P�:F��� ���c ��G�$� �!��F���=-�5�:��n��A����&��0��,�����>b��s�3���D�!�-&2R�Ág`��%�!T��ind�����Ýka�*�G0��	�U���� a+��N���Ύ�mD#	�*��䉚S�<��B�!�3F}�q���y������p�TF:�����u�N
�B�&�[A�
'U\��2�*{�$�e��������j񎀅M&7��n?[Q�c�p��~:�~n��U�;�q�����'�G���2c��g�?o�X�Aפ�?�[��W�!ȼ�ًkLI*��lݛ��A=��z|��ܔKM7F,�#*��1qcb=�.��ÄDr:�a��>�1١�N���ω��Ճ�L��Y���r��M���!	TU����߸�K��j,�E��9�k�y|A��~PFBΤp?�%ΐ�HC���@��A�}�,��O{6�no�Y�O��)�zF/�d���;���$�Q���d�(-��{z:#k�VxLz��u�HI�K�� �z��J ��\�ϕ��E�nY�t,+\G�cq�F` �.\({/<Zrh0�u��&�H����)C}�G�&s�k�oy;��MM![[̭?ݕ���P�':@㷱��neP ��1*�-�۱}�_~����5naaq4�X�Vٖe"���Q9@�C�
#����8��p2��qY%o��_��Ϯ��ޒ�J������C��5������Ǥ���we���*����Tk�Gc�*�CR����|1�6j�K��&p�7�%h�<�y�̒�+"h���t�|�ke��'^^�!���b��+�x-���r�Ν�Wn@�Cm�p����۶84�^��zw�S�[��̴z�&9v<9`P�����Rؙ�nv��O�����W�B�=�4{�c^��y��gU֙�8��1��y��#J���w�Pլ�h��C'�=�����l�#�u,b�kJr�o�����A�� �֍ז:�[ZzW���3҉�YQ��o��C�!Q�k���~�po�1��|�V#aZPP �qv�����yҍc�~��[^fQ��y\����ů� ~�JPT�3G�0-���H��Y��+%ջq��i��M����]����5����$:0�;k;�ʠ%�������}!�����kwr���m�H�|:�m~���������p�c�̱�w�L�Ҍr����?d\�I*��L������N5'�����MJbq�s��4
�_jT���٦�f������!|���iF����ͷ��D�����D�ND�cSC9OM���	���2�)��]���M�F�Q�d�:��xh���M�+]��9u��`����0]�|�5y�z��� ��bþ�L&�'"nפ�V�d�K�,�MK�m�����D�R���z�ӰI�u�1_}�<;<DHh9�D��x��F�E|�7�k.�ÉrN!�$�X�oQi,j�8x�D��L�g��z0�Ơ��婊4�t�*������Is�ψ�x����E�[Sc 	Cb��������SB�o�`}�J>y�;K�~��\젠Z��AppH:�B�2����*��5�I��K3Z�UnN�?(1��5���,T��aa I�KB�/�UiY����Y �ف)�r�m�b�	��J�`�H�k��߷y=�V��@���=���/�aoY���
Tۥf�w$��.qi�B�Vؕ��R��f�oT����O_|!㦓b�a��=׆�Q>��*��[/���:�ͭ�-y��F���^�5=���M[��@; 7W�X8E���_����I%=��?(��zg7���{Ԧ )�	!��Ǐ�DC��[	�/�,��yt�v��'���5hBlg�����ŖA=!�/��ě� W�E�N�	$��}t�~UY��0o�}aaf�P�j��^�:B�:��rѥ5�/��줎����
_���E�l �G;,��XD�E�W;�
xp�(_3�i�-G�	$�hN�Q� D)���
6-SAw;����� ������Cs�VD�v~~/��})�8���`���贬�{>��5�כ�i���U*P�{�'Y�تI���*�S�$%�^~�/��G�F�G���GӶ�3/����]E#c����Bqݶ���g\R���~_C�;��Υ���`_ A�#w���۸�\C���%X�8_���J���廄@m�#�S�v�q�k@%��RkB\|�{�Q�u,��d˻�>ʍ����7;�
����$��_CauC��m����qE����Jl��լls.����+O�Mۗ6� �@	UtI�L�|� ���BE�P.Ο_�����N8�Q���Ӡl����-�z$?o�Q�ӣEk=�R��x���>;�)~�<~yYzGD�i��>�8J2���w�j?�=��P�q��4;G�M�޹��� �K;�� �m����	��b# ��=N7f�Qr������K �l��~D����_��.Eǅa��c� t_�5�	��x1>}4�[Q	�f�YS��1�v���+�"|�2��)V�
dbq����ؽ��+����uz��v�uُ�z��=��@A���9�����G�S�^�:��[&�H����oCC���c�s2hGy[g�ֶz�����2�(ih��w'�}c��e�3���nv���s܄e .CM�@�4����&]���0�e�6O�=���*����F���ßG��66���U��C#�aЙn}��k,�o�F�ݺJu9"7���]���M��C&@�KGL^ "�uv���d'�9�%&*�N�M����fY}�+�(���8Y�����n��R�X\��V�CCL�Z�~��L��KaӼ�e��g���I�O����
�ZE�'�R�h��,`5RS��*�M�����;@� �VaP<a���[qq$i��u���7O/~���d9�zbM)�&]�Iͤ{�qz/fP�^8\xs֛�ށ���nm���Je|��h�(AI�ʔ�0��ݬ���`#$C�Q�~B�y|<`�!?�xTT0�Z�{23&#N,���ϲR.��( ;�\6��3=�]���~��A�X��=D���Ό�CA���C[D��,�<���S�����.�E�9 ���������u�r�~_\)�ʀ�= �lx���1�_#S[�~�0�|�C��H�����z�?bQ߶�W2m5�nK�{u��.�j����|���.��ʎ<�A!<402�O��آ�����V]v<���O��*���PS��]��ςE{r��[
u'KJ!ם� � x ��Y�<���i<����낄��g��A;�{�G��@UG����;nK޲�d�ֻ4e@z��Wҳ�-���k����D݊�,2����0�/�h�%N2�4k��~g�&����~���v�[��� ��<4tttJ0�F#�,�HYT�W+x�WalPkpo�Ъ����Q��f�x5�f�Sj,��c�eBŵ��"F����&C{S�K��,E��8�ךu��5�4x>k����:�v��K���k_���rc�e0K�ed��w�9Xrt_\�ow���-Y"r�rݞ�]�#�(�y
w=gޣ-
�S@|�hJ�j:�������ꀐ������.\��q�����Ş��+�YΟ}���QlR6��󪣎b�5C�Ǻ����2����z�ed=��4�c�˒yi�M�G��R�g�m_���pI�^1�'���S��^�U^��.s�7�"N)D�j
���
�yr�$�^�L��g�BaD�y,�O����y�d5�f$�RR�̑���<�f�:��C^�V\��0���!��1�Tϻ!�5a�~�I�wM@�G��_M���4��-Й�=
�������7�м�ޫ��!���n����xD�8����=;[��B�?�����'(�b��������
��-.��žL�h�"�Z䰿���d�~�Qkk5�E�|%�v���n�D5��ߋ���\�ݟQ�r
`H3Vof�>O�H����ä�B�I6��]����ژ�mž�Zh��i%� 2Ұy���7��?��͋|��2���e���FX7V�S��oy1���N��s�ԯ8AV�n����4�o�9�BF�9�o�|./���:��z�	<��=3z���|S��hN�����Q�Vm����`U�FHo�U��M��O���	=CC$�:]�*u�D{k;���cJZV�tӘX��U�-�TQSb�	�,4�aa6fۂ7H�=�L5��4�y�t����IVGW�͛�c=(��u�] �иIL6U""ǝ�@�ӭ6���j,2"]����'b��Y��gi�����^�`���-cf�����ɐ��[�d����XN��K�&��F�y��D��[��F�Ai��c��@��`{�DV�{ש
@.�߷x�������Y�M�*�:��/��Kq��@�Wi��^Be�L\jV�WQ�?9�̡�@V�,�ݸo���!�p����'����#^��m�
Y�'Ԉb��0������dOY��x]˚�f8��'.�����.�٥���[����w�M��\���X�A@YgO����,�ʨ�R�tqsE7نC��� �r�xu��5O�s�`�nI�<�l"Y�! ]�"w��������9z'�cQ0/PQ��_��l;��o�q�I��
e�H�/+ǻ����c�p4�lwT+��\�E�W�j)�ظI�nN�Tkm��o����v�އ�m6j�KG�S�g��.��3���T��>���A�y
?���Ϫ0�TC؟�D6<voOEC� j&��`T�ɏu#�29�ؔF��W���/�����_��/�'2���i��?���m�G9�I�.%&�#�7���Q�I�� �c��]B]�[L�6�g�F��-2+u�����z��I_4�1�t樛�R�?Z���2������A�PY�1*�W�{`�Uj^<ꮤt�a��j2ZD���`P�x6
�8ܡY��'��m��6�C���V	X� ��yb�	S C,/᣻�Ӯ��YB��ܪWB��Y��g��V�]�Z�1HU�.5��)z�3�I�r6�]���,���l�aH�R���o��}��n�ph��������L���}�`����Ȥ�-b�j-��w�yX�cM�@R�%� �F�6�,9��)�|�lt�"J;��w�qz	�Z�.��V+5�)�(�`Q����q��7�NI'1���$1�C>ZN�����]�������	
ӊm�{����E�!���g�i��,��\�X�X�l���Pk{�"��i������!��nP��}\���������M��+��S4p=r�c�7����A���7�;'����T���q�!�!�E�L'&���'�&�7b���=��� ���r�"(��;'MkF��i��;�~W�o�,���gQ��S�Hn����M.H,/T?��"���gf�S������v�%��y��J�}z�NU{��K>d��!�ݾ�O����7)]]��L���$OU���[~��C�b��r�Ƅ�f9.��˧:)/���"+K�wR\U=.{��>�&h�F�`�m��{������<��z=0�Z|w�)��s=����G����-���6 �<҄���@����E�R�<����B��W��Qr���K�C�N-��ېe챾)����������k%�Xi/u�T]��O0�_eU��+o�ZqM0�=�z�>��ș�-k:��T9,��R��
���uZ�.�l�:u%U��
Bu��>�<K�pU]�#�S��o7�|�f�S�os���b}�3����~xeT�7D��j�Y} �>#|${޾{g ѕ����IA[�/bT����ڸ��j�յ9�����N�,(gL��w�o8�/������'	����pX�F˛
0�N<�ϰ�N�/K�����;:���o�����-u�MJj�:
�}'��M����`�^�n��Aw�P?KFb�d��8��)�����6��z��~����bfn�8���<� ��&�A��DJ��[4�o��y�6�R�� s�����<�ʷ��]��s$a�S����㍕L�7pm��ɛ�C��ٻ$L-,�D��*O?3��Ԇ����� sq��9&&D{F��w[&�I���3;�g@���.1T���V��}�����h���Sa}�楅1�������ENw��|<]��Q�7L��
AJ�=�ب[�(qO�4�ʋ9\�Z1���r=&�C��/�$N�IΦn��.p��ڱ�*=��w �#�oX1Tc����a�b�՝��C|afS�St:d�-+q�0�o��;-�{�2o�Ov���T���j��Uƿ�5愷�T0+��4�0���Q��/���S�d��;�����[������g��`o��d�Z����n��k�s��i��]����s�n���,�i?M���E�_��=P�OFA�2�P>�ԍ���<m�gd�e�6��ࣽomZk��~W�[]\��{���d�OJ��?�Z|�_뮉��ά��<E��r��{�7����{o�B���K�]z��53��wnݸa0˽+�|g[�sc|�����x��M[�����z.��=άx��ue@�9�/{T���
��k5Em�9E�$b0_���� Z��Y|��2/P����xb,�T@�;[���K]���zi.ΟGZ���<�:F08%8���׺Ό�6�6��T[!�E��/�u*Q��aM���%�6�I��1qӾp~�fS�����/�����H7O|��P�P6���l�Gn���2����E����凧V&S���?%�E��:up��<{��bj������U��%�D�ƍFn�br�l��]�c���[�W��L�eA�L�v���|���;�ګ�:P�����-e�a�0^+_� <����m�r�ù���U6���I�K����U��Q'X12��p��M]�6lQѴ}�0ҝ����]>�FQ1�8����B�4=Y��p~⇊ aPl���o/�e�>g.��_�e�7�rW��n�Mh=#�<)%{6�M�G����D��&h��gs��3�_��(_�^��&�:;0]��mR$x��Ҳ��?j��;�t��?[��Y�4�<0:�L�Ϳ�V��VG->^.�P�H"GE���z����շC��l�p��xJ<@ԝT���w��Sb�W��<I�;<��ň��o���δ�SХM ��k�	��<��:)~��^Z���nK���;ik�
0�7)Y��2�6�J������X��{��2Չ��W�C�utMS�����׹�����o��Y�s��u.p�7"��5R~���k�k.��{w.;,t�OQ��C��5��ѷhxȃJ;8��MNjq�4K5Ť)��̚�=�T��N�w��vF�~X\Ժ�~23mX
��(�L*���-���N���˝S*6q��|������Ȋ�pj-g#��<�q��C	��glP:3魽���w���<�{L���I��{V��?G�O����k�$
0��>sI��1�ʭ�6.�- �s{k?��������y��	�?��#���S�H�]�ަ��P�y6���ϫ``�p��T�c���M!\5#Ęн.e}�|���MH"�t�ğTq(ú��7�.~&6*��4[�Q{pS���]]H]R&���5��kΩc�^���� �}���c��m+Ҟ��������&�b+�m9	��:3��"���X����(	����]S�! ŀ��Q�IOf*=�0��<�}��_u�v"A���L9�5���5�J�	����}�#����& uT����Uؔ֡�ݔcm��\-��p(0���
-�����Rw������%�D��^��y���skZj�t��*�VM�0�8�k	�Ev�RY�C�t�YQp|܎���	6n���l�{��Z�W~��xX��ҳ�}�ze�t�������3�T�O���>N)��'�Ⱗ%9�@���|���4�ũ�N��eVn��UqG�����`|�;�XdLL�>�.�c��*O�r�����<��\�qm��&�
T�t�!Q�8]6Ä4$�Ph\�V�J�>�S��|z0���E�v�r/l�`���o�=� ��bnN|	��ϧ(z�~�2��'	�h���VhH�����^7��B �bP����I�b����+�9�[w�8��7�(��iyg�N*��U\ƚ�'Mi�ʲ�̸����	S�Ǚ,i�laq�%%�-�
_񌲕� �%[_�K���g�Zv���=d
b������y ��%AA:����U���ޕ���umN��N)zZ���^Q-b�����<�Uj֣!��iUUMG� �5ϡ�Y�Xb��H��T�|����~?�?���+�˵�~�Z������_�x5��{Q�S轳����Te�s����gʳ;�@�u�J��\��V�Jx��՚?S<캕�ԙ���UW�/��y;�cOE�t�3���h��U��.~m�ɧ�s�HIYN|h�y_ވ��<�����Р��2+��.�|l+��Ess��6j���M��*�5�z�%e�6��j v$B�[&	c�K�i~0�6n]埠k�	�3�)1��Z$� ]��p���f(����U��A��uri�P�m'�LRy�����Jd7.?��������L��୨��̀�F��c�~�r4¾!�h���|Zl�.	0�Ý�O@rҰos!l�����~���cQ�^�ͮEG�(	�
E��v{n��2�C�M��|��D_���TG�?�F<4��ws v[��2�4�G�,��KHg�m�~o��$J5��Ԛ4 �el�*s�Ǆ��A�$�}|��Nk�~�vҀK�F�؈8��	�����;E���Į�F������݅��X��u��gyJl_�S2���"�Y�R>�#p������#O�;��	p@&+H��ܴ��&�/�����_�ƿ��b�4�w=��Xzc��V��E�k��P2�d��*��A[N�%��Lx��ô܏+���{�$��2���>�������^�p �;�p(g=�����Y���/ ��P.7A$�[���17bQc��9��ףۗ3�h���?cQ�T~7	ʲ����t�0jf[7�����@k�px�N����M��]-��~0?���lCQ�D�����4�S ��Y6u
�f܀��Q\n�Ex�?������v}gj�X|Nt��ޡY����t��6�2�D�ԞT)�&b*"��}�n��*w�L°4�b9���IW�Y��������	pE=�F&����ҋ6	��D��vW{�)5{<ڠ�P������tR�����7wH�P�/����yj�*���Z�#>�LV�j�:��L�������k�'z{�D��3R�$B0�Ğ?��Oh�ع�G����f��9ێ&����V׶����U�MY`�nO�u�*���Uwܾ�^�/��z�?�f�����P{{��ftF��:��"��mԺatY7d.,��u�Q5�G�{�m9A�H}iJ��*޽{���U&?��>��3Z��c�鹋Ρ�v9LwֶU5	e[���(T^p�ߵ�=���z?�B���\<[�!*�P�
�e+K4� �(�|;2'#�>�:"_VS�+3rr�ij?�{}�]q��3~j؟�R9\f�x�]��^�X5ѩ#�H&�\�Y��F��:υI&{�>؛�\��ý?�<�$-���v�N׺�nXF-�Z��J�(X���B$P;�ؔ��!OV�K05��U��7��.�#���w�An��l>f[����`7��Qr#��S�T)z]'t:@�q��<߲�L:ֳ�f���pℂ.0<�}~�+�[TN��I����5l�>e����K�sؿm�;�H� � �����k��ײ��`����)���*d�9;���k��NI�������o.%�~$����|�,���i�7kcnp��=���pڬ>�K��]�%uwM���8��7�{L�鬃4&��t�������bԈ}F��>���Å ƠC�ހx(�䴃��T��1Uq�O� 5j]v;�\v4{��υ���6z���\��蚕�jZ�����O�����p�St=�\.���3�e�?͠���V�<	�����H��-	 �*��F�Ei����\�s�����4SA�3�>��@LL����*g��V1 �+��0#p�K��鉷���~��b5��薿�x.�Ɋ��P!3��U#��π����+��~=?u9�W�����F���u�ȑ�B��BD_<�!1v��>^�63xn䌌]M;��?���,��wd�Q��T�G�z�s��٨~�(M��'�XUP@,�S>�z0g"}d5um���[��E	���6�;�[�5ׂ��A=9X��n�v1��Z�w��{I�˗�>>�^��K_-6��Ȋ�S���Qq�-��G�f��F2l�砿*��HS>)��nOLd�"��a�LV���B�"��q"D<[�8������K�Y�\�.S4���ϧ�8��������e�lҸ~�Aljj����lm�\dro}JI��y�u�l���T�sE..��=�7���h�p؏�����_��������!-��P�W�|#����(��#~ma�bksu�-�*��Ϧ�v~��c�n�y��l&eɕ3<8�d��u����U��.���-�SY��:NQO������ztkPݸ��;\A:��s<�u*�BF��������zt������ݸjd�Sߐ���bqR��Ѽ��?�pV6�5��mߡ�P��}e)�T]^�5�t���z�EG�c�zo�	q�F7��Ҝ�,_�Z��z�z��
�<�� ��[�j ���b~\�6���ٯ���L,^���'����ʣ��{p��k��B�w��bc�j��D}�fRBG�	�-b?XC�6�~���z�Z��$���p���I�O��w�/.~z�k6#��@=
q��%k�ujo��E&E.>���2����Ȧ2w��=3qIb?}5$�╊����<ݾ��׭=�2���A)�n�CX���ʦG%���J�\ǟr�T��8�+���O���&چ߻W��ʣPd�ћ�ҞDP��z��⋵S�dP�R3��Z6���σ��ܼ�[�Ql����*��׌� �_^�쐾�nˆ�i��s��FуX�#L�u�����#B����n�4� �C�*�����u/ߓ�MHQ:�"�%ST�����Cn���
H�Vv���!�����viq9*QM]����{e��g��u�O\�a*"x�@�m@����(��O�y)j��ϛ��9���������X�E��h�Du��gY���;|%�����2���� ��0/���_O�Ӏ�Y�]<��=$u��ҦB��cvg��a��]u�NS�z�|����4�4��&��Q�̜%� ��MZJC��0�!���$��k1���0װt6��)�ݽg�Gժ>%)����y�֪��EE�`�M�y�t�4�m�y"T���#��'����BE���X��9��O'�h�%���a�x��ߞ:d�@���D�����8&���{�ѶA5�N
v�w�;7~j�fթ Pk7�L!+m�#v�I�q*	�ҴO	��o�C�uKjFu���� P�^�qʷ/�����t����3�p|�2�}��R澸�)2�|�����D]���k�x�LN@𨸸8���U�wZ�F�})K�w�S�������-�mr����*G Q�3!��k?���-����'�K�������i�`b� ����B}��y��5
��B͝砆ⵐ*Z�g�޸����%ƀN9&����_��<X7�9r��h�p�/5�F<-n]Z�;`樠�����g{p[{��g{qF|ж�꿰`%Q��Urr+S{Օ�b�D�$�m��b_��x�lJ�p� -�g|s��6 K�������d@;�Z���m�.��FI�n[�vMO�@�7(�0�퐔�S_�5�/���ڶ��^
ǘ���S�>*H���czG��VgW���
�_�*1��ɕ6�����k�~���nJ��M���A�z��F�_�������6���;a��h���M<;'��8�-��*Hp�3R�������L�\�?���0)�F�h-�~�l��"���Qi�N�8pS���62�;۰�&f��f�:_�$�G�����^YZL]���ݧ����t"h����Phm1��5��q�Bd5��h���^ wTZ����*���"���n��g�e��ʡ�	j�bbJS���\>_/��ڹ�۪fJŰ�a�Z�ǇF���%�������:��~q�X���L1�W�u���z�j�-��yǹ�>k����y�B҇sSk�d�o'��Z�,߶�������!�(�-�bdu�@��8���.�m<���D��t�M��ϴ4�J��Y�?g��{Z���8^�Z��ŀ'�y� ���$����z�?oi��̳�}�	:m��/o�e�gN�܃�t\K@\�/5���z`� ���{�[��I7S���͍�7�z��i���,z��\��gh��+�`m�u|М|e�l"�A��S���LK^_�Ϩ���U���\�m�f��a��]�_.qk�]	WK�7�=ó���Эa��UuFk�e4�e^u���1�ה�C	�0�kq��(I�5ЩJ5*�,��5E�$@Y��c)r�vWW��F^���fA������l�~0-P�@�w�=,"G/n���۱���U�ٚq�4
���]����ܐr�<����e)PP_����伱�@�FW��V�/Cű��7's�o�����I_Nb�Z�a�Ag�:oO�T^��Jd�Z��-��׮�o���x�	eu���O;\������а�;�e�F�}�ͤ�0�'�
c0{Ԉu��^�����9�����'����ah�'���V�sr�%6m*\c��e��P���E�C ���H\ y1�</�>>���nwɌ�#8镙���X��ݴ�~�����B��2���A�f%#���\X7�z��Û�]���;.{U���Ӈ���t��E1���;�ce����Y*���&���UH r�RX�[��U�3�q:W�sq�π5���a�V--����l��(�\Z���:v��m�T�#�Ϧ�h���6F����������l��B?�ك�H+u煸����ΪTx{���*�=�O9.wQK�^~ ��q�E�K�d��-s��6޶G�0GU���y{�o���]�_��O_9����G�=�L�^�j����'e~��>�V�'�9�~�}�.��N��UӥE[z��?*�h8��f���������F�9ȟyoZ����c�ѳ�Ř٣/K475�1z�+�"��D��-m���F��#t��vuAH���{���� N�� �����'�n�1w�9�P¯���8�Q��[��?�W��*�_�����S�au�|˛��6���*U�e{���[��'��7����˨���|%�T��5b>�z�T/�JdL�I2[¬*�m��1���QyȢ��cz������As��Ж�ۺ����מ:���aO�9���
1VBf?۾���{�\��|��xy��*q�\m�@q��ʕN��Pm�>7���~�F�[�T��z������'`;J+I%u���Ee]�d7�\�+��&4}U��}?�+"����15��w��m�Ъ��ԝ.7�{�ű>{s��� .�=�Q��h��́������BnN���܋�U����m����[-V��=Tg`p����^9����E�9{�&�bjC����l��҅��Z^�'���ڒR	��"�Fj��o������f�%?����#��Y\��{�Exw�2�ѵT8�E���SP�ٕ�PK��8`�WoZZ:!5+����x���S����	I�U��>~��C	t�N���X�8,��T]��@m��j{1�E�z0�gy�W�%5�{Da���
!sW�^8���׋�O�П�r1�}�c��"�������������O/�b��ۯ��_�������E���_�v��w���w������*z
uF�A� ���7�;���'����?|;��<�V����K7�PK   ,V�X&�n�-u  #u  /   images/294439aa-ec9f-4672-895d-838110657847.png @㿉PNG

   IHDR   ^   �   [�7@   	pHYs  �  ��+  t�IDATx��i�eו��>���5qI�)�����Zjɲ�n�q�vv0`�F�8@~�W �� ��@ ���;Bl�c��lY�Vkh��5Q�X��*���;�ag}�Z��[Ū"�������ޫ{�=w��^��.�w�ߑ�w	�;t�.����%���������?!��܋?!���������f)�K�ҍX��$�f��aW��ti��������eZ��h��m�Pѥā���4�>B�"F�;��	]=���w$M�y-�16�w~O�����}3d'!�<}_RJ�!P��شꤿ�,;麮�$���^�R����x��<��/,�!�o��cS�s,�3Yv"��p���������g�ﵾW��]��|������ZF(�;���_�����voؼ��'����<��^�xS�����:����m=oT��zۮW15���?��O�/��G>��{��]��R
��|��yp4�ԬGd����Lp�LP^J�U����2OJ�j�Z���ܕw[���%N)�a�M�OU��wR����r��V�=�q7���^`c�B�u�-�e���E�UK�1�N��t<AY������?O��Pw�L��Z7��J��?��O������؇_xO��fJ;%�?�u{>���R<�*)�[�U##]�|�}Aɪ�X�:�(��0�T)�-u���H+e�FbYIݶRT����\T�^պQ��+{�R�s��N��b�ڵ��Yא*$�õ�_(*}n��f�w'c}n��Z*�M��4:�AQr���
����\��(d�X�`�=��jy,{{{�&�S��hC{n2B��~�?�߽��?�_��?�G����p��C�"�\K��_�ڏ|�K_=�T�*�p��AEj/�+I:��I�Q+�+p��WNQ:�J�g��@�Sq�;#�Z	�7X^u��!'eҶQ^�h*X��ަ�k���X�F�&���Iǅq��V��D��e�L�s]Le�(z�é��W���!sp�A����p���\�ZuG#PM�Q�BJ���d������?����������,���#O<��E���	�yp-�X�p���7.�&��+�I�9a���:���N��AcO��rp����:ڲ�{��X�zS_����u�S�G�h�D��c��C��(%�M?��.�%D5�s*��.�b��F|�J�Y��5�˅
���u�A��U����ua�������Q��T��
�`��*���K]���MƲ:�*�=p]�̟솃Nvv�<�ȩ��'��?��&��7>�{���b�����B����I3:�*�����R'�ꕜ��WK��3��Vܢx�:��`:�W`{��K�!J	Q�x6;��Ɉܵ�I��j0U10 �g3��N�}��J��8�b����#ٛ��m���RU�p2���U�RNw%NZS�JP<{X��jiu7�tqֺ+[}/��H�[��ѱ�t\A����9���nԅ�rWE���jmI�dн��ލ��L�3���^�*G?5��;ҝ:k�Qֺ5�:���j�(�Z�b�b���\��3O��~�S2���� 0�=��o�/��W�{Z�������z���S�ě�|����}�'����:�����ȯ|�k�Ra��	/���mQ	�ЫBŇ.�O~��ȃ��r��8���ي�������k�+�(
׺��x�VE�B��خ���;������s��1Tqb&2����/��\x�2��L��X��Qؑ3e��꼹ңU����]�U�����ʟ�����^�x�g��S����V�\�h�������d����}��?%�#�M`��u�S��_��Wd�� k�����X�܊�tUt���'��B���u��y��|�+kG�~_iַ��P/����b-���yLfǍ�'%mݵ>��?'����@5AJ8%R�J8$]U������O<+O?y�*��~��L䗿���Z��SR��c�FE��.��\߇���E�Ͱ���庫�������O�����:Գ&TS�I-�N��T�$��:�� r��z���P&�\�*U�+ǫҫ��Q٨� �����o���"��\v����oQeլaK���ve�JXp5c9V�^�J[wʸR����������7���Te��nqM�����d1pfT�^E+�F}��;R�N��j��@��x_v���7��u)'���t��C[�h�{B�{��[h<(�wKx\��qX�붛�؍nǵn�b�#�N@_P�<�a�����;
:%Z�_(Q[K�����Jf�R�Q��@	�O,�B]��M��B?�&���ٿ��U>)g���E�2����u����Qί��׋����ִ<u�J����	S�J^	Y@q�+Uؓ*ȴ4�Qk��t��2֕��XԎU�V�5�7�_��M�����9�,��0��r�ݍ���jtn*;<����6��t]] �vQ9x12W.�|��jjI������T�UcYB'胋rQ�x*W����ZjԮ�ܬu⥚���tc}�~��ʽ*�'J�5LX��P~귫�[r���V*~�c] ��n�1��8W�%�܎>�*S�C�;X�:�k`�" "�`��*JcՉE������+��*��lt��𮤽'��.4E(�0U�w�Ϫ�r�N&�J��:Pͺ���\y�ڀeQ�9P�:�9+�4��DS��xA���qQe�XwDQ�(��v��@�j����-��F	�r5�r��B�t�����7�~Kk�Vg����i%��6�Q�AF}v��pW?[_�>*S�B�V���Jm��Z�R*1�ӧ��kWTt�z����mT�AOM�b�=_����W�1nZ�m�I�"�u���ʉ�0�EP����F�&�|W���������K����ȇ?�����E�����<C��NH�S�S��+�f*�I���wdq�|����٧�������\��_Um��f2�u1Q��2S;|�� ,�P�U������C���:}N���,�o.���k�2쩘��\Ad�T0Є@��+��%y��T>��O�U4�_��_�׮�uհ*4����5��s�=��X8�26�PW���3�{��Y3
�6`�T�=����[a��,G�W�����/</���<���k�ߔ��gA�\���{��4V�1�}���%�(�cj��_�%��o]Qw��䃟��|��W���׿(��������{�*��ܴ`z����ۯ��|�� ~���}��s�\�����j��2���\\M�1-�CKS�W��/~�W�a5'?��SY?���_�W�$����ϫ��;=RDB��8e��ӝ��^ Ϫ�P}X���UW�ԍ*�F��X��]��;{k�*��״�0�pB�+�J�{���u��j~�}@e�H#35�hS���L��o�*��SSwE&j֭���������??~�A�/�,t�;Cʾ���!�F-�������U?�����rq<����:�3C%���cU�A�1%����E<��wO���JEҹ�r��Y���t|�!�|����չv��a/��./`�A�ρ>�X=cP l�3<��Bew[U�N�������sO������8�h��N���d�RI�6��ܮ|��H�(<�?)�9Rք�>Pm��T%U��(��!�ѩ����j6����Ͽ|QzX���D��2�Y@��,mf�qq����Te����i�$T���)���>�A��st��60��`Z�8
,
SQ���.(���޼�;[����?tS�;��pX3��P��yaV'������to|O�d����ړ��A[���!���Q����2�᧰�Z+�,V3��4ׁ�j���-��J"=���q]�
Q���,�L�NTfF���HE��[˷��	�� b����������RY�h��4Q��pt����G�=������M+p��Tdo�b	ܓC-��K�0G��[��7��F���h�O'N�11יLm�1�?Pn/ʍ�EY(3"� �3���u�4ÁjX7j)J�f]szO.�n��ĭʆv�Jm䑊���w���Hmp�X*���t��*&�&��J�����J�!LI5;�rl�F�y$KXQʭ�+��*W�9��~�Muؒ��C8c�{b"V4_�hOVj��BLw�r||��椇��ZU�xA� B�O0�PF�>S�5R_�`6�RO*F^u �CZZC��}��DV��
�xkD��f��p|]�/�n�Z*Gb+�r�wƶma�����}�p����eO9&D�~[]�6UA 3�.���������1�ա����J(5\A�M�C$3���i�bL^��YJ����	6>4&P/��j����@��Q^W.��^�����(|�Ce��LT��؈�¯����1��0'�)��{�!�|u����a���%�߼'D**�u[�x�I����|��VBN��c�{`�C������jw���������=y1��ĲM�)���	�|��	��l9Iйӝ�F�@1��E[�����l���1�r1�|M	�.p����I�%�&.[��U1"�?���ˏF.��[l�9g�'΄^�b��7�
}����(��lċ�=�'���aĒ��H��_����8:=:���n�pt#=�<vX�a�a-G�Lt������I(Υ�3��J�JE�q�ql?\k��@�8��Tz����-i�υ������g!/]'��V���<�ם��=>0�![�F˯�����s�����)����)X��)�.�a6��+q��m� /��HXp=�
���Y	]�e�뙉�$�hk�8�¸���?&G����K~F��o��+R��}����Cp��6��r�&c;f����8����+�t�ӊ��pr�Ȝ%[p�׃�Ֆ
*QɈM�7���8>8P"��gY�����[��I��Y�|/���u!�����2���%��]�+�o3P^�m��³@Y�A1��ǒ�oІ{�ޱ����y�@h����v�?��n�HN���|� �k�q=IA`D�����i����	F�J��D%�cj��!�᷉�m�������|��V��r�Fr�O0�]��P�J}3�(wzv��r�o�`��� o3�$s���B����n1�1,��>���K[�ol�q�+�~,)/~^H�s:��d���M�'�����n�Cp�U�+���5�讒��D͘��Eo�����R!���FS�\w5�l�"hr��XyYr`�%@/�Vn˂�x��I��i-�Ct��%�A��0�f(��߁lX���$KpZ���f�`]�mȔU���#��X���A:��	�!!#$$p<T��"��&2a
�eh��}�HsR;���������`�T&����kP �L���F�$�8��Z��@*�����Gȅ`�֬,VpI*�B"AAޢ�4�N'd�
#8�ǎY���؜N]p`{R�L��`���dpzU�
�%D�bg���&-I=0�4ͪf�Ɔ��S}���n8̡�5�C��XKw�yw��w
���@#��$��}bf��>@x/�ˣ�.�ʵu�Ơ�A�ԑ��H�G��H�u�F�����ಋ�aa�V;��pgB�b~Gj ���2UI�5���U����lmQ)���e=�ٸ�|�L��{�}tW-e�􉮓0����,��+t(n�0G�n�6B�C9���h9E�HE�ޞ�Z��? ��mx��ֵ4��tJ�`9	bA�s:��(AR���{*��,ή��B�>���h1^|�
'|���&���K��f�b�d�r��y�w��QQ��].�2ra�� vyrsRܠ�x8������{�/�C]w;P�&"/�� �5@J:�aD��=��k�~�R��@��6����1֨��6�k~�QP"������a����P�~�$B��	��{Ő�D�+0i�W�9ww����������< (@SN�NNHx���m;3: 3�� �3
�u�δ�!�d%n�76����Ǡ@1q��J���vP���P6#klb����sr,�ХG��#��&��T����>,8�������Sk�1Q�vq5�oc��L�� H&�{��+���֚���<�U��f�uƐ���<K�~�����]�AC�[6��Ҫ� \�F���9F+&đV��|�0nb� ��6������''s�Z(Hd�c�Qۘ{���mK%U�g������.��L�@K�i"���ν|wpOJ�U�J�"$�s{Y�ъ{���lz�0#;��`,>�-NFD��h�4��ᖉX/kd����ԢN��u��zv���[���aV,��#,\YXD4���Z�oN�c�!J
�z�@�)��G邇Q �m�}���ݮ������e)&P`� &qf��@>��th�3U���.����0�-�+��
8XjS�3Ue�c��܎�M�䀦"Kd��M w��.A~�,��Z��0W���"a ��l�} o��F��>~�9bu�I�)D-��z�M:壻S��v|�(�U���jz��v(����\zp�"#Y�i� r�1G ��z�h:�%Qj	�9�F'G��r#a�*��#>ʰL��Ȭ*|nH�S/(C`A �;c&��h�(Ԗ^s5�s,>ŋ"	<��Ň(S�=Nc�T����Ȍ�������J�0�t}�ƥd|zO���� N���@.B15H��U8��b䌒3�Q��J��2�������ۥ�3���@��ݤ���YA�r	��r'���R2Hr� JӁ��4Qg��M&;�0��#z_5��pj�O�6&΢QMԝz!ce�f\�I,��a�ߓ�Õ�,�AY��	��
+�B4�R���H3���jCƋ��_���0��#��3yM�4 b�P<��� $`�a�к��\U��˝GS��qx��p�9a�f,tfU�<7��d)�?;�M�;��!uU�����b�Q���+���D��hK���
��\�v�q�6VY�8K!}^��a�1H�t��@���= RHn'7�ĈGv�IV(����W�޶#�|Ki�bI���$���]w/�����tb5�4bL�ʔ?�.��d�}�1P�\�t4��b�V�C�kVy�����c�����N��� �OK�3r�Õ���@0[�Y��V���D-Jle�˝���@������V�QzS/x���f9�<�eum�䖏�c��0��h��\���5W��*�Dn7QX
��~��q۸0�)'?�_��&�Z�bO���3k���>��-�`g���'��;�g �Z��Z��ڭE�,�DA�n��֢E(�/V&��<�����cg�S��Xpш�9ä�!���xa�)���d�"���X�l$��Q$VV��@����r���`�E�"L���%�Vډa�	u�ͬg�n��G���Li��0�|1iJ�Ո\8�'���a#.�}/�m:j|v�kT�bwn��O�0qb�>.4�ض��\oKx˹�H��A�S|s,)`�k��h�)�j"��<,�of*;WK17��β@!�����̾���T�b�hfz���;�	0Ya���Z��
u��ˣB�1?<b\>����Ib+j"7�,3baE�T�v�=1R:�m1�Ep9VU���t/��	�LLo�y�',:;y�9�c2X�9P�����踕�ru}8��x��R�%�`�@�N*YO&��b�� ���`+s�bpXX����4���=H�z���fT��w�=�ݝZ�۠t6fȖX�z���ܛ�L7ݤv]�x�y�oZO�0q[\?��9/���sJ��1��S�R���>c�-z��.<\���	�����хAu��w0���QQMXgKj�����9�l�PT�����#���]R�wZ'�a�+��ޞ
���&�i�x2��Gɖh{�%{�w�1NJ�G�D�24g��K�,
��I�v�g;Y��3;k[+���E����p_h���;a���#B��mhN��DZ�2u�J1ڹ��9l��R!l^����a�%ND�����Ќ�%�3ci���G�yXULV��h)���@����߄�%@��eTߋ}�.>�G=��	�G $��s!��\���:�
}��̑h���-�ROw�GpQ��-�� �N���	�k#���r���|s+Â|6AX37	��1���ڪ\����q�t�8=uȴ1�F��7�,��9 2yE	���u�т�Of1e���	�߄��8B�nE��z�56:t�{	�{�,2nmse3����]����Y���U�,��u,�@��i�F]R
�O>�9tט<�Шha�d��{�,�P8KW��O��}8{3�ۯ��n9�����d�'��Ž��cٚD�pP��zɢ�JM?�΁�o.�f����H/4�F'x�Z&�W�B�Du�v?�`RZV���ؐ�e��	�t�� <�͸,�����!��M��s�6,�\S
w�8�"��`�dA�K� Y�>"��� ��x<V�ʌXȖv~;�g�,�V�¡�>����,�9R«�@��*	��&��#���.Nu�)Z4��c��BÍ8�X���3+s�6�On��$������F�/9�yC�v`f$e/q���}[�=B����d���,�?A�R�{Ö^���B��$T�/k�^���IT�DU���F�������� '̖(��6��U��$��Lv�Gg�d#r
���v�{ZC'�G�y��2�o��B��	�&�T]'�5��$.��9r2p�C����˦6i2�?�vx����^����(e�{�#����s�y�q�����d�㒈��:�B�1� �fᒋ(�2l�"�cM�g]k���:��,Jx2�wM��E�0s����e���0�Ye�|��[��|r�cI��SU�L��pe��׻�0��3��#׋��G������:�[�n��y��Q_�b5b�����*��*���	��}w�8���p؊��k��������V��lp�}��߲�gqGl�<^ߵن�b����H_^�<�$�S(}���q���2qlN����[,��8��]]��N�L(zH�Υ�S[?2;�T�~,��{��I���3���>Xq˛�(c��?m��e�X��D[VKj��󯡪n���9�u�%N���Ot�4�-Vp.1l�E��R��Dw���N۰� �egM����2��9�1�K�)�P^����m\�����zº"��S��Unc�蘐e�\Iՙ�]�Y���;E��a�-�N�($�7B��d�'Q ���q�K�	��Z��х~e?3�g� %ژc��7ߞ��&��b��F��:Z�\;��St0��~��V���X�ƌ.�ҙ"k���-K��M6�?�P�Q��l�e.��B�L\��új���oD"Ϡ���s���JF�u.�++%�9� ��h���U#���G�e��W 8d�~kz����x/�ɢ2�?������C�(�T,�����[v��P���to�X����T.�o�/�[n\��A����P�41�A$A�|)�C�ܯ��tA���=p�Id�V@�-��0E_�#��+^邟�ϝ9�JX���J&�1��9s�-x�a�J72S�/G2B�����+�NJx3�"�4t�Qj`��oK�m���斣�o�ܚi7���t 4»�>o@�9����/����/3n�	+���@=\X�p�@�<�f�MK�~� ����I#�O��A��M`1�j�0t6��	E#����8A?5�yM�����d�;�a�b���&S�۱��
�f��ypa��.�N0/Ъ�+�%� d�]$8�	t��5�)B��+Ƚ >�1�Uwf�8h���eaT2	�z�)x	�xE���h-S7F4̩T���j�ɴe$���;��*��	�u}cowj*�5l�����l���s�N�OG��2����#���ј2�y���ã�X�C�`���l�N�x,	Vjd	�����{]�a�k�2 �t՘��x|�{@!� X`T4��r l��'
�����sb ( n���0A���w��p벐���<���xT���oJ>-9p����y)���7�a� ׶�iWt[z;��mWS��kF�w��\8�,��,׋߁�R:�$j��t��`������E
�p���<��LB*X�?_�׽Q#�[h�PV;��%��� F̞48�ʳ�Vk�X�~=bh���G���J��Aa�7�k_ a�O@Kh�G똔�М��Q��jv��2 ��x"����ղ����ǞU��2;� ���Q��w��NfN�l�8G�a��Įy���}ۄ��[ V�X�}e4���D�h@���N�0*��7q{�͔�Xk�h��H�\�4���Z�3�;B܅J���:p�Q�B	H���{��rr^ȵ���r'�s�A��6�����R��QOߣa��j���W�6�m^4�A��tÒ����Vb�tf��w%��T)�����A*f��)�]��<U+s����Q�J����01�'�У7�;@i���a�v�2i�3��g�M.�^*�$�h�������Ȩ�����Fmv��a��2<l��6ұxGЎ����e�tK�iYR�.���#�=Ũb��]=aˎG���J
�!�u'D]B)�!|���h�X6��7.����(]���ø"���%��2�����*�Q��EƎ��o�Ü�����(@��(F���3hT�0AW��U�T��_Y��^���z'(�l�؀�^;`
jI=����w�qg;��7��"Y�b�r���2��Q��h�?ϸ�k�a#����w��*=b9l��"pl����e��B�u�41��s��.��Y��B���$-*1��G7���@�e%��_��+TSd ����$ngӀh0��R._q����0��$�R�@Q[�.mp�x�!C��1.��=TK��dk��+�P�ˀvш+l�
�ebg��-<�m�$@�W)3�l�8g���.B�96A~O8[�,�����gl��K��}r�߳�Xr2*X�C��5��8rk�Y��x}U�d=g�`=,��esN��-6��J	�n�W�M�v��}�4���ܓ��t�3��]�0�"���nG�B�ַTY�q��V��a�@��`�1$���~@������B`�x�G�l3.0��,�B2T�{�.S�1�M���%X�K<�jܖ�J���XE_`M��	�d�k�Sbv��.��
���neU�F�������.ae:LpG8���˃i���C?x:9��gX0C��3��6���"����?҇-`���~W��%��b���E(F��h�EgX�jU��#͊�N�V���e�b��B����W׭ܶ}���)��a��������ż���J���>s��Wli��?0���xn�`�o�{�����eJ�\C8:u-9��L�2a��
�|�x��L��l&���Kff衑�!���Rr��[/Y\?r��bf�]��@�y�h�GR.�,ʤh���v|�ǒSAd��I���w��+Ļ=�"�g� �J;+�a��5��7UL��dc}	��Lc%|Yr�wA�r�Σ��,-��GM�Y��:����o�رi���8u�[�����G<3"��g����d���zf��O��څ�`�7�__E�S<1�Jy�Mܚ����h�>8��c-�gE�fc�����r�|�b�k�v(����q8B��ĺ&�q��\�6I��	���H��T��z�rNQ���vY���E�R�g��=3Wά�AD����.AɎ��X�%�����B4�PƓ���1�\��9�c�3���(���*��NB�X��.��(�@� �Z��!x9��t�b��l�f��he��� �P���g��f/r1Q�y���òb�X��B��q;z�[���X-Ӆ�,ܬ��,R�Ʋ"�KUǄ
�w (�r̒�����yX�����2�0�V6�u�{`��	>��~�d��Ea�vqt3��ɂ��xl9,�(�� �"�$���i��	���F��Z�5U�@��0K�9)�$��޸��΀���J�Ύ����ɲS"�̦r���Q�x0-��R5-����`�K^�q��j��	(�i�f2~�_惶ȑ�B��oJO>�ɄfvP+����.ͪI��$��錴�Гm���䛊��[��[��"��ڭ�.|�Yx�u^n)��(�*��+#
ۥm�hl���w�!&�����ʇ����x�w��|1&	�]��Nt4�D{�����~�0 '�J?Y��*.g��K�U��̲6�!�0�dA�a��v�"�!"~�}_1����)���y���L�DY;
���_ܺS�br߾*9+�Cp��۩�^G�B:x��ob$N�P�I��X��� �O�-��e�yr ���i&2�<8��`wjI��<L���@��!=�\�)^����Έ��r���8��j9��?93�*U��X�&��&G��B7x�T��ĭ / f�#�ES˪��+�î ˁ�>��v��d�����;T���Cȿ��0yv\����2����� {N�Q,���HA�
��
��\��^an�0Le�ˊ�g*E��E�	�(�����H-�b��h����ӣ�>*贱`�mخ�B�|�X�cDe�f8D`)FhF�-`e+5Kw8c'���h��pG�`H��S����/��ְ�=���%|�|�y�M�̰�dDg����o|,V��
>�4nP.����X��e��2��z��6��_��k�-O�o�(�qӊeU/���w�bz�s���lW,͵��]����=rc	�
�nB����������$��;���60�"��%�� 2MG�4SO�Tq0�wV�<�vM��Ɋdr��		����bZ&
�n�		���o�ڭ�V�$��r[;r�M�Y�h��K�yWc"-�+2��v��	cEx���q �İ���yMq¤]�Az�������(.j���R�o:�Ln5�*(���jt؁�i�����U��A��ћ�� ���Y�#���q<"��|-�S�+�ܶDz����]�E��W����)�ά#m���C����"Ӗ\��m��4�OӮΒ����-Z���]�e�܋��qp��o �pM̥��#x�IB�C��P��C�*�r�"94�f�El���6�79v�҅�Ky��75VV�g��Z:���׭��&���&����!���ˎ��Y�>�wrQ��,�����Q���b�l��I���(x���Ak�H�Eg�]X���4B2%IdV���IF
94��}-LLGb��� RR����H�`� �f���2Q���%�W�;���^Tm_ᤝV2Ȯ�v�[�V)Z�~m�8��\�����JnT\��	<�<W���Y��V9�l�:bH�w�����5|(��_�_'k��\�}:�xG�&N��13��
y��d�q���bȐq1�;���2�]a<��}�K������z�ԣ�,θ
�Y�|6���Le���k�_�ŉ*��X&�.�Νs8��A���be��:�VB�j(թ]ZY9���R�����d�3��EP��DF��g�l��Q��bzӷ�����_�M'5ԝ��ER%�
��:�=�۾4_E��a��H��x%r�XU�z�k=4 ���ݎ������!�L?�X�J���:��匭[�.�_�V�@�hu����8-�ޔju�C�X��]���.���-V�iQ��-�8�����~�٘3O&�L�n� w�[o�
� �m�cJq,�L�~b��h:�\]��<>�*2��x�ag�.�ǉ9����ú��y���h�N�wґ�d�΂�ڰ�I9���d~q�4�[f}�m�6n����$�U�ա�q[[�'��}#ά�V�ӹ-_��>@+-j�nإ5��齃�4�`�P�u�J�0#<��Y%�Z�	2�)jk�a�1?�����L�Gh�_q�U�9<�"��Б\�M1ԅ�.�Z͡`OCg_$z�5�����@xP�2�B�vjo��̿XD��+9�*���ῖ��sB,��-q��7�����Dy�Ie�'FMF7m6=t����*��`�M�
*��a_6����]ʖ�[udn��-I���Mr9#��daηH�܉.����+�J;��9ږXȐ�U�IwJ\^gEE�fc�4���(�?�(X�ѭ��!���ʹ4��E��l�ׁ������&r��w�3���^�lF�f���zG�jrN�-o &��ګ �ǌ��ݐ�(������~V�����Zw���\enD����C��Dx;r4�<T��B�N�@��WW�DìJ�D)빶�S���C����d@�鵷��}*N�e���\d��Y��6�Xv�;e�����P�����bc`UJo",RhU����xW�dB���J�q�8g��q��^2�]�\��ԔeA����E';��-&�6hJi�3���m��pO3]䭂���)�tө�]��~P>�i��]F�
9s�;U�Fd:N�.
��|D.�T�F(�1������\�4<S�=Q+T�ȣj`U$��&�呼(6U��"��"1l��[sN����KXx��>oy�[�l"����-E�l[x�RSZ�\�kv-ȩ[u�=��t���>�Bd����u�L5L��yR�`H�fDv����l,-\�\�4�q��a.p|&�47�C�	ɻ��{9�2��N�W,ۍv�Z$�Ds *{wV),e_�+��mѲ1��膇8w�y��9!v^ag�AP�ۉ�2X�1'�3�3k���p�`ֶ��D�#N�Fq�0�D5���1h{�s�E��V!�C�ܻ��(������.�S�բ19k��� C�e�{�k8?�"Db�л63��c��n�Z�[�[ݵ���݈�-�j�)"�ٺIF�D�{����B��N����L軉�;utz���'���m�Y��������Q8q$#�����""ٮ�n���qR�$�T��C�&��[GL 7k�����m�	��Dr,�,���_[��ޔkz_`��ם.j�dS՟<�f�PdPj���D�N
)�7-lЙ�ø�B���L�h+[�`�>,��i��i1�h(c�.�~��b���|��9y/9�M���~O<�3���M���5��=x)Z"�Ȱʎ�K5=����|)~ �'ѭCj����M���U��΂��+[)��P����O��A�e��vS�s����R��{����8��L#����cX��̢�٤�*@p��z�� ��z���ɘv�2ؙ�`X�9W;�H�?���֩	mY1�>���St�2�';�č��N;W�L�7Ȇ0��g�}
o��6�;y��^����Gy���޾�<]���=���D����<V�P�	(Y�w��tx�+��l�����#�<p%��dmDuJ�dʍ��N[�ŤI �mv�����9� �^���nN(j�|G܎+��nx��V�������#*WI&eɾH����(�Df�������k�� �BD}����W�ƅr��hz��Hm��~J��-V��=���W�[�8.�#*���ᄢ�h�R����%��7��V�$��[�b�v�5��~�oY�\Xv �&��]�S[?�L��B�)�hE0l{���@��ꯨ c��'����w��7,�/X��qW�JL�V�8���ؖ}��W>���t����s]�b����v�s�k�p܉�n;�s$ B���Z$�P��<�["0h���>f�cE���yپ\2���&�i@� ���O������_�#���]α�ޒ�<�ΠC�����ݔC����T(��j#{c��?1�u��P2�&9Y�ؙ��R��4{��<�е�_��.�Lkck�mU�T�7G�|Kş���r�=�����'�@����%��z�����q1�cJ�O}�����[td��#�V�vc,�ɔ�Ȉ�!��>�Bb���@������A�q�X��f�`2r��jp<� ��1��2H���m��"T̘�iß��]�����9��������\��%��l�dIͤ������5>��p�{�1����u�G�5��#�O@x\ʥ)opu��<���N4@��x�0� ����L�k�]�N'�53��v��	ָ�s�0w�+�.�� �̀�f`<?t��6/�M�G
|�lz2I��dX�,7��[�^`��`.�6�����!vw������m���,h�ab:9�#���9��2�<��är�/��VV�C�x��M�C���"@�d�%�s�*�^��u�H0��։�>�<E���Ax��=lZ�9lNOF����D6/�H�I����rҽ+6����C���wo,�Σ@�4�ͦ\}˨0����"9� Z����/�L�E���� ����cW�����Kn��cn�Z�"�ɚC$�A�w���f�l"̮!��tژ�v[��؅k�K�o��d�O@��F�Iz佢�d����(X�\[�Ε�&k��Y��"J섙�h�N��Z��z%�6�lW��+�M,��"��VN^S�[�%8�4	�;�'� �	�M��Mض1v,�n�WEmG�a��*��3my��P�:Ή2��U+5
����.u��&��k�IU72R�q�D�c%�PKa��P'қ]�V]�:1��1@�,�5
��āo���ȇ���"�{�O��Xe�p�@0��;�@�����߭�G|���Q���]�Z�n8.�LM-�uc�0��m�����=��Ӓ����*c���:�k�|���wCx��b��JdW�����K}�a�wp}�g&��b����f���v�d�S�iBOI8O(T����b���r��	�!ܣ��@��|!˃ci�IZH8S
%2�	��\�|U�ျ xIx�ƥŚ�k:�.�Uu �~]��B���oV� ��Ѝ[;���mk��z5�^����#�p�0k�Q��w<���U�o(��!B�#��-����\�6\��`
����v��ߏ�P���?n�[u�c5@':Ik�'%�2Z;A��2���}�@)G[0�1�ɓ���֚1ԅ�8�����mW/AԬ]t��7���й',vD�I	O[8�J%�Գ<����
�Yu�x�:��+R1���+��P*9.�N&"�p���j��֠`uwY���`]�fi�14�ѿ���0�Td�7�`��v�S��*��c��/s�^b+�7|���V��'#k����$Z7�}Ψ��Jʢ,O��8_�k��e%LQ�2\�d�T�⨄�3�=�ſ!|�r?/+3�P���%��i��$b�e��u˖�ּ�
���>1zn�[S[g�ά�ܦ��㜷S� h��*�:ݦЁ$uο5��}�aP��(c�x1�G��Ѣ�^�ݣA���k؉��J��s6�vt��z������'���]����'��{抖�N�5����+k���T��4��q�hL�ZVX7�)J﹙�&�2���d��]f\���-��y���-;5!>����C2N��Iҭ�Z.b��8�4׬4,Q�Ү/rۨ����	�����6�yz��g��ڼް��fHs�.Ő|��m'#��89G'9�#v�^�*���p��Z���/s74�f�����HӰцl�`�Q2�%�`{As�� �yEۚCU��]O}����aQu1ډ��m蠰�ۄ�v�Vn⟓ȹ�����a�"l�}ͥ�&g;����Քm���<|�}r��9펙"Dt�hv,�o�՛7�����[z��v��M?���ț:�'g�v�U��"���i��E�e�,z�Ƣ!���R�j��LƷֳ�m�B�Xl-QZ@2��E�qY�([@���2��l��3)�M5o����F}xM����<,��A9�� X�m����SCy��GeV?(��y]^���\�r]�����Έ㔫���D,6��z�S�6Z=y�&Y=z�ĺ���!���u�:�Vg��(XL��έƙI��J��1b�Pz,"VSTlY�^+��JR섁C�AF*��򖧔� �z%�NMe~��7)�G?��<��i��rj���/�{ge��.���z�M�`f���rz�>yq2��rI����Fw��d���ʐ\�XO#븃M�~�Z����#�j[�Ě���j+�v�Ӛ۹N���w�W�:.Y�)o���?���L��L���Q��Z�q(+ג��7ԙYUC�Ը����Se|I1c��u�,o�ٽ�|����Y%����#���O|���O�):1�V�z]�ׯ]�/��o�|���}�	B���M58������]
/؎�NV"�r}���K4L5k�5�}���iK<����[��N���wO��+�)��4n�T*G��ӋC�ouS�.˙�\�uT�0d���)Q/����S���iY�㕟�I�D������&���o����K}�������g���?*���G����~|�u+QF*J8�'���N�7��=y��<���Py�ڥ�$�!7Jڲm��L߄�څ8����J���Y�+���P�ϓ��~�Hn��n	ߖ�-^Z�JR�e�_��b��uy�芼vY�-dG��1vC�n�N�P��f���\��oĉ�G�ЦϠ��;7Y�����+����������H>����՚D��Tj�a���,���O�^�w_�G<'��s�q�,����V��0v�n�j�Λ!��#���1�!�����cluS�ʗ�	�d�Bn_�5jrN��k��壋krvyC�Z�]J�y�ّ�Nx*#U����b�zu���X
��eeg��VT���=*���2-�*^>,ݷV�
��%U��\��MX���ާ"陧������Z@oޜ[���xD�\����|�I�=Ҏ~��Ys��rt�������'�Cl�ؾ����}�^���7�jq<�D�[X��d	�����K��Rf�T^����T������t�y, ��=��}�U�.����Sc�r���*�[tOBC7q#�kU�ν���#O?./�YNM�rn���r{�f>+�K�{�V��I;E��CF����?'���lG{���*����5� �����Œ]���#��]�3*VS�>�2v�5��������%vd-�y`q,��CUƧ�X-����;��� �*���Hv'8�b&�S��*p�����9Ƣ0���%��П�1L�=�7��ّ쫒f\>���c;`֓��
�x�e��NM�����C�wT��2�������;�}Y���v��8"����iyw����6����r议�)%j�����;�l��4�V-%�d廢��`��8����������x�PM��@k=��Xlo#���D}6�` �'!ptw����Ǧ�b���Z���8~Ӆ9���{dq|U���oȥ�Z`����⫯�O�b��`Q��:��S2��^�O�����N�gHy������[�N��'�l�*�7��R��e%6�G����L�S24N�1��%�gJ�n8�q���|�8$``�>�.����J��X�N��y�=����AW��Wa@���H�����d��̡*顬�)�������6:�[�}�{����pd�>��/N�9�
rU��Y��f���81H_V��
Y��x#	�V�ن`N,C;ZX��Rf���&%��� (�bd�p0nUz��+��C�7?���vy0�\}��.�N/cG����5�2�2��dﴷ;:����ysH�NS���b�v\}k�^׽EMWX����d@��j�6���fT=á�X�is�2䨜������tS/���E�X��2��Y�99o>_���L<u���ƛ�~�T��pX�PQ��F�-*�8OH��/�.G�H)��54�F���7���X�V�t���\��z�5t��Z�^���g2Њ�ڪ a8��d���2�l�3W�휖�r.St�f��*:-I�Sn��k�=ym�/���ZsnM�>1�M	�#�~�?REэ��N�A���5��?���6�R��(J���q:���r!ce��/�*�u'��s�h��^�
::���9L��L�goWy@ T��ǽ�m��nh���h{�~5E��%��תPU�\P��7��!Z �v�!�+�LTV��9#�<}�|g�\��ʑ�Ȇ@(L�rH���-����ɣ��Wo��7oȃ��<����xP���]������?��f�Z4������Z.^�(��ղ�g���֍\֍��;+�MǨ�ݥ�8k
��
5�\�tc���n�����Nš�.,�V��AH M�L$r�;�:��=Q���oT#��J�s���)]�	��(��w�b��$p��cZ�s\�~(/�t^����K�廣R�����%������m�9=/�����o����I.]���.�����T���t
�ϯ)��MG�ޛeC$`lbAi��c�:�� �-�+s�n���Ȱ�qΨ")Q3S�YM��u$Gꬼ�3U�(b;Ki��!����X�O�䪊�U�mGa1x�Uy@j�o�)LG@i^��&�~v'���,G�����~�1�ݝ=��E��k����;/��9Xv2�]�^���rniݵ����x��4�<i�&�*��8�8+u�%��<ua%��fz�ž�
�{;P1ƕe�<�E_�+/�Կ/�&�� �  D�B]�y��e9f��N���>��ف(��(�>C��?[ȿ��s�~@Ə=(�/\����<���d��C��@Օ+��P���B�5@�;��$����V��[--�2,�>���Jn�b�DfC0J�C��̨�R�d'K�C�v�����u��m�{N��ݣ���9�m�q6�t�hU�.C�
���6��l��&�ɭ��F>��Y�$��hĸ�JM=�h���`��J��Ǌ�H���[�W����v�M���ԺQ���7����X�=�f_�v��o�7���\[�rШ�G<�r�ƣJ<�:��/#�8����{��F�R�"��<�BU����_F�m�y1���T^>n�X�&�_x������V�iǧ�j����Y���z������<&�1J�a�^�CU�+:(���8�&#����F����X�vF�廯_�7�U�|�!9{z_
Uԃ�>O��|�������p�K�*��ឬQƃ���Co���J��S�TMb����؞1BI��Y-���g��_��N�W���,嗾�=��ﾩ��`�!qK����?'"�lv�[5��z�F��h��1�H��̎����豣�{�*�C}��`���a0a�a�S����= ��T.]y]n��}�f|�P �X��옋>�찂���lƄ8�I��Jul�.����f�~�U�kS��u7�/W��8ݸ�r�����L��vsJo��Ԍ1��ポ/�����<G�xH-^��1+��L	2��i*�D��r�V'i.��7݌rjoW�a}?�� xD���ҕ��9��a�~r���j)�T���p�Kd�TwJ���c�������!��C�.,��Cuh��VH�����g��]��l�T.\]�'0��6_�~�܎������e[,Cj���h|�'x���U�ݔ�r>w��*�������am�F�o�H�nD��)����9�*���g�vwd�{�fb�C��4�C��x6j� c�X?�o�Og��3���kQ�X�7<B�]=t\�{j\��k�б-h�/P���&�Y+���v�����>�V�����A����ngDmnq��U�|�6;>��s;j"Ѫ����b���o^��w�)�1Ӏ�[bw-uJ��O0W.�b�*� N����[(�jdV��rA���Z�g"�^����P����6;<�"b��Vɩ}���7�d kJv�)ke���K˻���g������d�Er�F���;����*H����'�/��3z]�zM�I-�z!g��(QU"���\^Pw0ڧ�;�ӟ��^�g\�W_}U�J��\�xQ>�̳�lw������b��ޔ��	-��Z3z����|���SO������O�c�=)_��eg��<��g��͛긽��8������J�ğ��2)��^�v�ʯ?�����Iӱ#�t���&e�
�������H��u=a�~'��[4/�v"A,_��]ʃJ����>U�y�7C>�#��G�Y��� �{�C��#�2�}������۸��׮�3zV����r|�M9T����?����l)���y��}�S�?���^�]</�/�y9\6���������xn�n�g?�	Yݔ�j���?�G�_���ď����~E�z�9��g~T��{�o~�KLr��//�b*�?�Q95�+'��KWԑj� n�6[��srw���s��>��j��(��?h�jF���,�y�{�u�v��{\�~���������E����d��\z��s?�s�S?��(w>(_��2D�����#���_��_���?�Ay��o��OX�i!���/�g?��ҿ�'������ܼ~ ��c���-)�.���|�O�·��7_;/�x�i��/��|��?��)��_�翡V+��N[w�V�Ҳ����)�ME���g����jZ�'��w����T�"'��n7mF�A�����2���v�����0��?����^�o���?�q����������a�.r)��P�|�j���'����z�If�Ν}���=��g�ܙ��s��>&�����P���r^~�gT~쓟��������ß��3�e2��5��x��I��V���TQ��p�������W�o
e���d0}\��85�����g�H�w�D���hP_�#ۥ��%Qe9=+��Uy⩏ȏ��?,/�q(׎����������gd�s�|�sP޼rC._=Ro���t_F�}����\�vhU�E����?(K�&�y妄��������7y����99u�=d��_�pA~���r����?xEv�{^���q�/ϝ��z���*�������_��|���`؎*�v����I���LtA�z�;�h�2�П?{'��߾��y�������0k0P��"�
8j��I\?Z�?���(�������/��5�e?��UV��Pa�r��y���s�H��E��?��n�yY��9C �x���ټ�����+��+�گ?/o\z�%��h;:���ã#�@F��/��|�׾Ά_�җ����̤����<��K򘊯�7��S�t�qT6��;���[��,Vs���Iԋ��=��a_������voߵoc�ZR؈_z1��GX�=f�do�'7���j���/��{CUd��1O���=x�Z�Ǉj{��U���!F?���r��i1Qb_������^M�W_��Ě��cO���7���N��>���U����gO��b&���9�߁^eC�M��_72@x��
g�[�.�>[�dto�\��_K��?���W�wp� .��e|!��G�7�̓�r�Ԯ^�&ו����3'2�%7G*3�*��c%zO��UVr�VMZϙo�B_�U5�ܶ��tF>oOEL�'�,��xCMĠϙ�G�ڵ7I��gU�TT���HE�Z5��ǲV��O�P��G�mq�PcA���O1��|�*f�����wJ�{<���*ض��Z��������J��߼fEe�]�*z���zv������g��}Rv꺫�������K�����ng�f��ae܌�~J9zS��G��x�~���K��\����fR�*-uw]|)Rl�y8����ꎰ������[p�z��]ݹ�H�d}��1�w��n�|q[���v�A�#KC.eIv��j�]~�Y]zE�P��0.j,�X�,ܪ�7�����\]�b_e)��^!��]��q��S�E�G(Z+b�5�4'�En�.7uw�Ï��u�v,���<�pe�ߧҴ�"�2��avK�x~-�����{�E�z���֪�n����C�ecxz���S5wB�*?���0HF��r&J���G�' 	��^�kUn���"Wt�TNV�L-n(Ӣ�]m$���CI$;g��B��b���'O<¿\S�qz��y�!ځ^����������<�E���4!O��� ��r���Ee{���j(+]�+�Ʋ����U����x9�ѯ�K��@g@�s���=/ŉ�d�VÕmW�:,I��ܲ$ٷ�)�����r[Z��T¦�x�_��k_%�>�Z����[�(�z�$~��C����ÿʒ(��{�ɍF�Hb�M��� ����<���9�5�-�N������}Nv����/]]�k���y�J����=�����@d�r���N:*D�;A䂸ET�K�U T� f�	m�x�|���gA5vb��G|E/�Y��U�����3�ʍr�8�<����\�|��k�㤮
~���Ɓ~'fI���F+C<}�_�{�����@��v��^��wF����l�ڑ�0+�?�dEd���<� �+��PZ[Y��Dhk���+��Kd!�Nԏ6�qu���l ����S�ډ��1M���Ί�ge ��H96���	%�ϰ��
 >���޵��u^��g�˜��s�=��61)6$M��Z���R�����_��4o$��<P�$����}#B�T4��N�_�:���ˌ�s9�}��g}k��̸�N�����h2�������k�o}k8�Ҁ��:F}`|~�(���VF��@QĹ_>{ݽl.��u���ok��]�w���"R�!��H�r#��R$t�n9�
]X�d��Q>BO��{�]��-%�%��(F*��M@x
A7It��-�h��)D�}������/�ǩ*��M5 ߗ��5�.�>\8_���/c2�al���P; -5��)A���9]��	�L(������Ǐ����|�́��[\;����џ�QD�=�횙�\���*�}�{�*@���R䚕3o��:IT�מ�85�l��S/эפ��!i��u�.w*t��7��R7�1Brk|���sV$+[��&wv���>�®��ߥ�e\;��}B���Aj+�(�U(�`j}A��JZ�o�#����O������u��R,�'�K�Bg�xzpB7+d�՚���~���/R��<�˗���cCT���H%�V��a,>1E���H��۷nѵ7����TU�G %	��.j~}�Vi�����>??�0�7GSt�����,�½W��Rq�=�M�,�w�V�%����R�T�K�"�+9�kl�~��*Ҡ'F���-���7]e# (j�۴��,��.�x+�[햦V����T����쫻5߼y�q� 7���T�U��af*P�C�Pg��L�	�U!�Vw<���%���yỻ�Ԉ�Y)�[�1D���t������ v�>�w1�.+Ͼ���J�+ש�mѠӖ��LK֮��xH����\�Em�N��o���+�3jq��J�'�(T�.|v�&M��A�^�N��cs��s ����,q���9�K��s��d�3% K5?e�e�&+89\��T�اj��D`FW����t�=�(!�$�K˹����!�l�D�u��	�H��qnu��Y��msT�7)�����8��'��A���s�����6���lҁ�io�:k|P�Z����n*P���P�\�0#m{eP8�z���Vg�Sf��o���Ǘ�eF?U^*��FG���"pT� �a.�/v+�5'〔ȉoq`wG4k�2mkM�C=�\����[�5~��?f�T�@�0��&���1�*�%c�٠N!o�5h����}���:�_�B�ܗ��[l�h��u�zT�kF��ݻ�q{P�B,��cI�/Ǳ�o�U���{��-^�E4�� �^P�ݔ�R�f1�°$T�XvEA��O����9����k���a!�%�j����HL�}P\�I+g��x}�4cop���ϡ�w3��п�(T�eڢOAL~cZ �hh�1�eǕ%P�W�.���ƞ���3�jx�g[��ԝ�2Y�]Y��bz��Of�>��T�6n\%�s��6�_z�s��|�	^YQ$�EΪ1����!�_�B�|�nm�3�0��	�����
�4�h�����t��+����� ѢM�`w�I.h8A�ϝ@�R�2��4�,<D��=��õ�Er���+��)�
�E6�PM��ܸq�+�X����s6�9�R�mC�>��e7h@w�������Zk�Dv��2E���6l,��hc�!~���gM������)��;O8U
6n����t@���8�)�Trmz�/t����ۜ���=���8���`�Z��M�C52�en��>F���o���k�����hbn�!dC��
'�`���"DbP&��M���㖭@H29y>�T\]����V����04�Zc�g�i5�d6Ne"���^�ϴ(TL�T���q^�Ż?D�F���8Br����V]���{�RD�A�",���)g�������-�M��5��I����p�V��k����UF.~��@֩û�T&h|� �ɍ��L3C䚻�p26�j�璁E�-+E/\��<��=WS��Z�~W�9��e��v~�Do Wzv P�^L�.�С�d[]��th�üXy��Ð����y���i̻���@���u�j�И�:	U��N� �F��gL�t��:���QW��;2t��H�ʁO5��n�w[ +*AS�p]҂��F�6E�'FUeY$�ʩݎ�@� f2���a��������{�@1HE��/kD��{i��nRXm�`D?H%= F����V���U=�xbx_�12�nN�����} 7ؔ2_�ςJ\�z%f�9�C�f{�*���H8���t��`=�	An���,�Ui,�H!k0H� �TMvQ���0L�h�yg���E~���K�INɠ�
���U�v��<���ӃY\EQ�OS!�L38BZ��Kkk�)s{Wï��[WWWV���9���<AG����.�c�T��QKyyȠ�X��r��ic��w.\���C�y��0}���TM��8vԇ9G���Q�#U�����_��J~H��دҮ�9�e�Zv��aB1
�2c.E�{�t�<ml�Q�Y�G�?BSӻ�,�k�������
M�ʁD6'���Θ_ZO��ٛ��qG(��qW�W/���"��7�Jm�|�[_<4�[�{�pjf�q�'&4]��z��c�l�J��cJ�?�[:�]���+:����/���6!���6�e4�`߂ 1��z�<%k��	[�#Gf��������W)E�M)P2zB��%M�}�e~�kT�]���)ZX���I	���^�H�O?T��Y��C!��dH�=�ǂ��F?��o��p�fۻ�҉�7N����o�r�w?�Ks�)�l�����itc�;��]�.4jh�ms�G�_#�hQ#��(k�7Z0.}� E3�q�� ���U�jrH6܄�tJ����@���G"�D�g:V�W���`���%�Gv8� م��A�¹���PY��Jy�j��`�����������/�x��s_{��0<��N�h�>���]��=�{�7��O�N��� \b���"h�F�BG[�tW�~7�l�M-��	���؞U~B>�؈�7)<�Ɍ�S�2�y�u�*y�1F;�(�1毲��s�#%G�V��M��ª��|����V3�/�|8F���k����_���$YۯD���**o�4�������e�A�|:!qɭ^g�핕s�/_y��~�<}�?F鏯��}v��g��x���n<Y�F�^��O��H��+(��/��qs��9EȎ=�T�L���џ9�SO>�t���s�02b��$�%��݆Y"���:o�42��$Ju|Ȣ�I*��uDW�����Ũ�Wr|l�ErF=���*� ������[o|�ԩ����z�k^��c�y�y^����c8�/��"E�%�s���W���K'>�Ч?}W��S����l�����c��݅f�W>�},@ �g43�d8n^�3��	��P���J:ZT.����]��'_�}�YB㘌�e<ak�﵉j�Jasԁ{i��N�ǔϳ�@�w��n��;o�$/��g�B���	M?�՘��?�Q|B�D�eȇdH �U�lK
ַs���3U��:����N��̠�Ky�}C�,�LJ����6~�:��x(�/�~�KEPb�tU�^ͤ�1������/��}�jvW4 S���~舆n���T��瑞eк/��=������	fvQS���Wc"�
?��l��C�m��O8�K^%�� ���&�����e^���?9�R�5��'���8M�y�:8�qFM��h h�
�H_"_�&f�_H��0�{s�ӷg������e ��@������Ϟu�Ï����o�8���=��H�f\%����v6;Q^�Q�s����QP�\J�K�{2:(���/­Q�c�9�Pp�8C��Q�z./�J�G��G�:q�."=9�D�ȑ�D�����Zj��%��E�U�\�S	L�ô@j8�#�D Z�iV`�/�3
���� y~��뾫(ȓ�$�s���?�kg|�ه��#|SQ\"�g�y�֠h������Y�Ҫ����1B�($�ǟa�^r�H~�O��M:��ٵ��\$Y�Y�t&�|�܎H#$�(�4]~����c����ӧ��C�,tvP{G�Ҙ��ƑR�]*Z�FʄX���bɮb\� ��A�M����2|�-��G]�ET�8�� ,�P*u\�=s+?�kgO����l�]d�lX4	�8e���,��ތ�˩���FZ�ǱK�Z�$�afs:J�7����l/?��Lʍ��wh��$�L�ϓa+�ʩ���1÷��+Irm*���]�3Ϟ�EqH��s"g>��9��PI����1��&�3�f��sG�KJ�2�!��5eM���^�)�7;/r����(�]^����'�;f�W���'.������G��azp��� O�x#œP���CH
"�5z@��������%!.)\���].+BR��ڕ�J�<r�Qͮ��8����`��[���3�<���Η��o�'�������8�٠���-����D�������Kg�o��Ǵ4�r���F綖h���,�ͨw$nPU^��N}��/����w�;fx\����,g'O��ş��3�y����澊�׭��F_RX� ��u[s���La����3�=ꩪ��M��3��\0�S~�l���+7��߿��^;��Kg����׎�'N�zai����k�n<]������5��q:9�����W�{3m��Q�9�����#S�� 	����A�ɜ"��JNZ��|p�����_��ѓ;��q���ZZ*��'|ݤ��_����c������Vsi��    IEND�B`�PK   6f�X�j�� 7q /   images/3afa6c98-60d7-4a37-9aec-be07fd386e0e.pngT|	8����R�$tN��J��%������&���-J�"KB�}(�JY��6c�!��G�I��g����*�5��y��~��}?zz[_���&&&6�׍��X?01�9||'�F_|:�����a�t����_�7-���>R��ku41�<�y�������=����%GW����������U&&!&��&���Kָ�ލ�)�N�>,ie�8z�ｰ�Q�>k���]��cr�c���e�kw1Cο�n�r�<��oL���G?[p��?t���7F��J ���}��)�u�������T���%�RtHQI�Ly��G"ovf�}��-��4(pTr�}�һYH�j$�A]�`��eE;�	��݅'�b%�ĦF�lt/�DP�����d�����sՍ�s���-�����/y �ȻX��e�g�П>�J��=H�m,T�k��kT]�t�K�H�`����k��R3�2�Y��O_�{��X��&�T���]U��+�^v�����sq0��96]�D�,潕�d ����6h�8��Z����-1�r���vsѱ��b0彄c�@��)��|�,Q����:��0�����o�t-O?�1�rͮĤ^h����#���M���@�g�p�F�(�J����pd��k=r��{ �zq��-MN[�]E�>Ò��!{��y,��3<��i8^j	G)�P���ʉ!!��[W�JՖ��N�����b���4|���N���.kK��t'w���$-���##��0ֽo��A�k��K�^/�u�w',T��}�E�	�i	��O� {���+m���.�����bmic��w��1��c+ۋay��؜=��H����:�޽[Y�^ȥ ����m�m�%{B��|F��=\��뚞vW[���.��h����?}n���ג+�KE��[l@ af� ��2_���X2�	�n����O�~����Ql���)v'A;1��7�}�Q&��&��#�d�^J�%�wxϩ�"Co���^3��ٮc�$�4b�K���#���e��ʴ�'z����f����7��f.o)��4�;�%]�'H��ĳXRˮ4�������3�q�H"��H�b�þ���BG����;���
��b(�}��De�0$��H��G��j �� ��C�*��X1��D�eE�@���]�,�m��*�$�QB�g�X�g@@���b�q����j�x�˂��ـM��BXep �r�t�ʉI���s�n6H��Xi�"I0��|,#�&��t4�/&wͲ��$�����Ǉ��T�iB�f)s����9�"��'����wB@#1�[�H�=�Ge���y���m��_7�:������ �����A�`a�O�eMS~����&��&^�N쀩ϻ�oʴ�D������$�(�Ѻ�CbC��<�t����G28�H䱹C�xK����� ��	���tw5��D�b<�ˏ����"_a�B� ��B��#�D����ŭ�~�~B�`�@|)�Y��r�L&gIϕw�57	��Z��(F��<W�g?�L���fz���؀g�]P�S��í"Fw�JLF%*R}ߤv�'��L@ri�%|\ǖ�pb�d$�i k�w1�T�Y*�,u*^��v����6C<	b0!ּ�"`K���7��C����Mlh$q��|�@�%6-"�k�OF�&�~�Mԙ]_�0Ҟ�Ԝձ�5���ќ���8vT��d��a%�8�r��3�N�Q\�Z�1:��N�䆸�B*�qx��P����t�@5?��_�0��*9�{R8�q�A����u��E�c�bJ��z�J��D�N�S.t����B�@�/�� �gh�[ [�H�����;R���So''�GqK[���51ӦT�/�����W�*4�k5���_a{H��^�(u��:!
-���Ƴ[
�,��Ä	�~X�aQu�~��p{<��S����*���詎?�A�-}ۯ4}	�S��bJq��pCLJLL�+)財E������[LA��VJ���D�Yb��������ހF{����A{d���������@������_��mQ�C�ԃ2$L��
�FZ��F���~M��q#�ā����׎�7�}�ۨ�ѕ�Q77�����mV�+�ҵqҡ����z��J�Oco�i\�ߐ��{�U�>�l��|��o��!t����������B8v "����>��jF��F]k�\�ʐf�c��1_����ٱ���K��I|���NG��1�JLn��/'�*�ˡ��5�-ڀ0r2={�,��)C����/$��v��^��������ׯ�n��x�����خ���kKۓ�N�Q͙�B��a�˟�CN>�z�Dlh\�C���nJ(Q��������6*:JNV�<g����5�Ԯ�x&�\� J�j�jltۿ��RS[�@"\k���+�Z�]i���GG��i�VG����s�V,a��F%�U˒0Bsl�!���U!;��Ш$����J����e��z�e'$�ܠP�U�Zo��jb��j�|��������9��N<#s������Yt�����B���҃Z�&�!,�(�<uj�c�8���b�ɦ���'���<:::87WXS#�@ԕ���/�?���N�����~jnǽX;f��}���	���Z�*	iދk�}��/w�r�T�����q�q%&JU/�M^��x��u�b\����QфYÄ����n���S鹈Y�Lmm-�P&+mث���x�-h�n/7%�!d(Og�q(v=��E��<AAL�ړ7�L/	v~`rw
~��ؽ
7ӵHaS-z���#�b�C�cw�%
�U�c���!����&�y EnH�GE�=�*�AA�^�sjR ��u\�0p��,E�b�v�-C���������������~�U��B���?ںfDd3��yz�*��k�QY��oPgnk�2o�	�)^k�f���:;�=�����?����	1�����];OI��5x\���������yډ��(�1ٶߔ:����,� �t�Q=|��ufu��a��]�L��/����jj9?~x�%�A��o�q�DL��=��Z�x_W�8'Q�2f	���`I��P����?��8����d#7�A�?nA �x�E���!el�%�4`/�����:�!���uZ���������ٶ�Д������D��z��g�4�l����q�Wf��?��bd�~�?؞�`��!;>В�l�1EX��`㤱��.pr>b�.�3ҵ�w�1���L^�e�h�t/�>����xezi8����KHioo��U�|09̤�T%>p�l�xk��S�#�ѣe�cɴ�6j�5+�����6k1��l!����D[�#+����=��O������C�Ш��}Lk��dMˆ�#�X���q��FN����9�Q��I���k-i�q$���1�s�q��%���2��\�6*�Z��.�%$@=�r޽����x��1_�@#�����..z�P! ��"�q,kD ��
���{��_�q_g�1�����S�@B����ܛ�Ǐ;�ʪ�Wt޸���!
ҧut(��9Kc8e7��3���Z)�f��;v��iK�{�4=�'zY����Kr��6��ntaI��c�y��?��Ib��acK�=z8��x/}^^^K+h��]S/S��7$��iIr�zE��5z����Ծ�h{���ݲZ�gDR��Ӹ1�?U33�3	����J����9���5���[��K$�Or����:�������Ȼ��H�U/�G�h'g�[ ��i�3�!,W�B�ϔ8�"�h4�=�y�c����o�)�F��fb r,��>��F�M�>�V�C�Ղ�"һ��؁��.�����8��9��h�hGק����9ɛ�2␋@�@��|\wղ�9ğH	1��l@e���Je��.~���{��)�2O;��x��n��9uXY����k��ɽ.���#��5�IW�+x!��,IP��߭׬�|�TC��~�-�а=�J/萭��7^�?^VF��F^Ώ�Y@9d@�S80�j[����̇�3H��mi*�Á�氄����/��k�t6�:¦+���k@q3����[R��:�����<=udd@�%I��ef�|DM�ۚ¹�R��TDSSȣ8���'��IR[��E�6�m����0M?����%�^�XX�#Lл<�ƔRP����O;8P��7��������m��t���w�l�^(��X�U�?)V.��@�U�c=ӊޛ��Г�I�e���m���:ꅎ�O����p�ף��*/�mi�tm�w���nsљ��OY�������x����F%��N�tw;� ��B��X8���>��K���j̵��M*Ss����+��%�.B*�3��	NM��E�C������|a������n�����m ߙ
��N���u�X�!ݒE��B���]����cZ1�=.1��jnW$�d�����[Ub��du/��(�"(Ky
�n�d8���ŏ?^���9���R-��fk:�q�Az1`3��6��L�Z��XrLa����r٫W����[� ��D��}}}n��Ds����k����R�4��vn��M>�<@}�6�4�"�~�'�z����/��OK��fwl[;G�X�H �"%5���@��K'q�*�z��K_��"�����3�+����N���*��Ռ�I����m���_��to���e;���M��
ViVV �.!110:��Hd��垆#��GC��X���X���^�/���O`2����Φ����*������D4�=��bDDc�-��ì��m����XjK�]i�}@\��=��O���S*�T-#Qu��(6��K����/ȩ_������Q�xߜ!KLbJ
bw���UW�
�����["��6[���x�!|�0gcs��@�/g���.)}��+^Xp��xbg3�9+�?��b[&&fy�r����9m�{刧�m�X�=���f�N������0����P=qw`�&�7S�GAyoO���9�FءBr#�	ai9*�PYY)86�>Y����N�q�]`���3�g)�c������x�n���R��PD��v��A���܁�>�UI	�� ̀,�Hl-{4|�(�c���lA�b���x�M�k�P������)H,,,�So���9�i�}����ـ
�C�g���a����E����vK�G���Ǿ�@�g�!��HW�R:�x7��� �R��sxb::������k�A�8�Z 
;,�ĂM		���_�/��5���i0�����UF6;�/���qAF����J�`H,TH7\�ۃ��d	�C���sU�T�Wj�R�(5�3d��g`p��c1�?Y�|}���E�@aF*j���NCخa;|r �DR���|.������"7�l]%����V3�l�]�M��\k�9��y�1��#���i)��j�%�\�Ç�pU�P��U0_׫�RW`U���#��{��M�FKWShC��f�H�x�_(Q#u�H�;��_~U�K���\" ���	eZ�\��c���0��ᶺ�3Z�����$:������8	T{�Jo��B��
��^����獋���Rrm�4M4S�h$A����
H�����/O4ѹ.:�����?�2�p��;'	+��@�~zU��5��~�r���#�.b'�A�j�>�>y�-����&^x�S*m�ɫ1�p(ۯ�2�l�3�q�o�Be�y�Q���2��ͩv���rpB�v�Y���[l'P��B�C>�{�St��.�-��!g�c�.	���!����73�OW�UlT���_��ڷ�G�ro���*�t�6V��p㳁�V�����-������_B^�MӬ��#�C#u"B�N-z�!�����w�[�0a�9t�r��l�RD��Pi����?|��g{\��WR$&7לJɣ�ベ~�D���\j��I�Ek�	�����FW����O�*⛮�nHnb��8���^��\J}��A�Cz�=q���	k�6��-x�#k[���MV~�F2��t�p��*>V�Ua4�ܮ���0-0���ߛ���ⳁf��0�p��6�mBl��q75c����M�V�o�X�v��hd@y^�U�;��)ymg��4g"m6��\���q4}u��\�V�Y:���l8q��򄲲rW$;��v1|���O"1���J(f;����ߙ�~6��E���ףX4K"��P���Ļ�d�ݫB��^؏��g�0���4a"1M�`{�`�qD5QO���:/����qqq')b]��u���H͉z�.��]�`o�-���ɲ�$�D��v��0�&O\�<K���FPc�G�C�bQY�e#u��Z�)�xq3�a�nue@<�>q$|�V�����]+-��W��a`���;*� ﶉ=��bY62b���geu���3̣�������+�ŋ�b/9WH��h��_���.�>�i�Z�brk�	{��qs%��3zz�;���˿�8} �d_�M4�����%
G� (���� L-��Ѷo���d��O5��b+�����I��֓�H��Q�B!��]�:1�ߟ����~o$�hs�͟uJ1�Yy&&Wr*Ի��Gr�f��D�Ի�:<����_�s�V��p^'�ב=rm3ǂ�cr	��{5o?�F�p�.r�R�@;YW�s[Wy#�T,}�x`��}*��%r�u����o�BWl}��+���%.y�;�ЫFE�;����N���>`7��z�B���K6���^t���y�Y��,i�s���w�r��A��I29dϖ�2'�50��P���< �$/��9F�xT&&�Y*��f�w(oa�' �oKL4z\���"�Y@C�����kmg��݉��:���bT��y�6X7�k���Vɋ�g�|~N{=�P�}f���Gc%q��@[[�+�C�U�k)�p�� �t���$��{7*1$�Q4��������x���+�|Pz\r�m*�>E>�w��X:�d�7i�3`�%�u�~�!k�^�Y7S7�RVL뒩��%�O~X2S �',Y��j1�*[`%��s�n]E}��5�pJ5��)��J��UBg�D�}q�gOA9��jp/���ID�r^<���F�H��l��'�r��+�&�RĿ�'dU�6&'��Y�\L>���NN��k�5�|�C#|��:�d�dP$1��L`~��<�Y��Q�e�NJ::�?y�U�ci>�<�N�u�tQ]c�l��§�3S��"����{��m�c>��ⓔwḑ��|��G�E�+Ĝ�l���(W��$�O��k��?�9:2��Ë�n��Q���!I���}~>'H:���URG[�\~�_�k�������!�	9.��XY= M	�!1y��x!T�L$7�����؛�>�%�k'&uc�����[%�K�~��ȑP�oT�H����1y����z�����'��eJ�4����Ѣ9��`w���7(�,��
��Y�)����k�Z����̍�-9�U����Hd���+�0 �#���`�0x�?k�4��.��I��u��e;}�d$=��u(��YZ@�_�{��kj�Y_9�� �?��o�D^�<J�V�s,v�l����I����Y�"p���u�G���_g�}��FA)�"p�Bi"�W��aX0P_>�����N}W0��kXrwT�)U��D �Ĵ�Ĥ��Gv����О�
��B:<<���kIz,��r����c錪��+��͆ʞ~��o�i4`S��~c�S�.�fj��^:�P<���<��pn[_k��|�U�K��:�(tؤ���b��	���D��p���{Z�p_��+��Q���Q���u�M�D�#��PW �Ĩ�w \V�D���� �c~\B�RA�R�J�YA
��E
�i�^y?d�⶯���A�oҏ�/�C ��.4c��JM�J_��-2�5&�S��T���퇿�ª84�=D_��ec+!�P#���;Os畁FMP�{�ʼ���hVE&���������+���FF��+�M�[�9��`�k6���cY���[�	�>n�c��G��}�ޘ�H![kW0���Oց/rNV�� )�����̐�֠}�*L_���?-���E�~������y�u5�Ǣ��$N��T���m©I�{K[�B��-0���/���{6����@��%�c�6bB�c���Q_�Y�{,���$��+u�gu<@�gǑ�Y�����c �V\c.��Z�7n���}G[�D�}Y	[�������|5�����Z[Ƌ�\E@}�IY�?@�}s��&F�#�r2�H�U��=!����z��򍓗<Eô�N�\�����.��"���Ȕ{�s��L(7�S���ؠ��?�Ϊ70=�u��#T��ЄWTp^���;��b����c�Y��-��	��̠���h�١-{$��KtS�Te���1��$
��:�"�%==l � �F)����J
}�b��_�]��z$�޷LG[��)�� ���{�Ѿ �����o�=N�b�. uۃ��O�k�Cpp'DiQV}���,����Μ	���PH^�G�e5���4N%&N�eY`�M�� ���8*�� ��'{�c�"��7p��$|ڸ&��2�C�C�l�G%��x\~'a& �ݓ c��ߛ�w�B>���x���bv�9��u�����;�^c$x�om�ɍ(?�5�5�@sUUUy�M��gD
���VZB�)���B4 .}���5�4g<�np@���α�@�7^�m������}��κʘD��2���+�u%�E2���A��bA�M���x&��2m�����A16�[P�����+;�]�Hu��u�}BK�t�9Zm5�$���<Q����@W ��_H�)N`���R�Q���	���A�!��f�/<�Ϥ��GEEɪ\�}�z���d�r�W��x]�ɬP^^8%��@��� ��_�| |�t��)�x�z,�^����,���~=�o8��H$Y�ښ�!H��ޕ���,3�~�(��#.>�r}���O�^�5ꗉ���Rfy����.V���p��k.@����γz�֝>Q��ת��jq�F�C�]1�IɅ�.�#�O��+��C�)ej��gR9���ҒS�/-u�;i>-W��[���~��m��
[��BR�ɨ)]�c���j?��N��/���<��Cl��L �����$~W�t�hеV0yc���,�`��i�� �y\4(����q^A<���᮪[WܰߞI�m��Mx�����S�z�Ma���n����<�h>Ax�٩m]�^΅�x!}��)������tB�>[��o���w�)�o+�l8�@^b����Y#��p8�8tŗ;J=S��C����e����Y9�R�>\���י^$'�S�n뀹Sz�nq%s���XW�S��x���(��|?Sc�V�i
����'�'��4����$|����giNO�-�e����f?b����� �=�q�V�����K�q �D�����!�§/��������g���:;|�^�r�p���d�#�2)|\ܪ?�k�p�0}�x�]���i+Pպa;�j�/�n��ST�q�u�iC����ދW��m<�S�8 ��b��ղ����=�I3���u��kYx'zk�#3.�u�E/S����Ew��xxy1�?�w��y9i��d���[e9�lV4����ւ�SMC���U�,�c	�`,!t�d�ᮧػa	�7�r�zU�vv��פ�������t�@��d	�Q��ge
37�d.&��:��GP�����_���������Y���E
���m�k�;�x�r'MS�kn�Qu��A��^�Ҡ��������_�׎��C�[�z43t׺�BeC�9�����yTܗf�ʱD���iy�qBxo-��{��M����+���(�W�M���FkW����Me�>��e.��1C� 3�#Z-�G�Xt2i�F�%C(!W�EX��#j������OK�ǒ?0�7t������H�Chm9bO7�^��
l���9��n&~�����Ŷ�_w=[T9_Rt��D��	�R^^�rQ2�X��c�E"S�d��_����w�r��r��9B�A��D����6�Ča@���"KE�=���F��0]F�,p�y��f���Eݛ����_1��c֏�" -�)ht���9���\X��e��w���Ӝ>������B�*S9p���
��.GL�<�@��=�ֱ�/ҏ2�DbB��n���V�Fd�������?��F�D-|�`q��x��c
���[ȃ2f�i��]ڗ6JNK�]�[|��viuB9pj��)88�21L|L���<U!C}U��Ω���~DI�
9�JZ敻�nk"?i�u�.�k��z�����^ʞ��l*�`�qm/��LK �����7�߄�?{�������������O;��b<����.?@ �^��P' k�ڹ�zF�4j��A4oЏ�t��RZW���!Сx���I�XЬ��,������K����ʆ�7zՋ�V;`{�A� �ݜl?R���H�_f����ـ�2�X�зH֓[��n��6��ϸn ��u��S0�c�WU0��)�n�'E,��]��]W�h��6�;�zh��dT�������,�C��e���lޑS7TBˈ�O�H�g(��j�r�d�?>����r���'���>&�Xi���ݱ@1���o��,*3�ѕl*���G��������p�{�Bd����5��9$	�|!s�u�VU�03�n��|�}�D�ggI�6�_��e���A=>	2���ze�g����ۤ͝����/rS�M��$���V]Y��;ԡviu�:M{^�k�Lc��a��d���1�ßΜ�A'���ڢ�{����$�hB�:�/u���@���� ��O�"}���ݤޒ��|�X��I�ORA敘k�t�^���V�Jo�t�$��Ҭl�L�bA�Jd?���5E�QH���:�����:�Ҝx ��s��øW��ᣔy!���{�U�h��\Z
�O�����OR�����h�,(p���v>S�O�����8z�pU�����hW����B��C9�"�I�w��3\W3��v[�Q���NM��yv���#:LC}�w��v�m��o8�bMB|��+\�e�̲�IS�?
�mZ�� vOf�&��Hj��-=G]���RQݣD�*v�]m�h;�]�IT�;�9�Jt}Lo~����Ӷ|n�z�Hjn��'�<���?�Z���*�wֱ�`����������s��i{�o���Q���9��>�Y$fe�v��������7�_��� *]kL���I_�mh~��k$nk�o��-���@r���o����z�����nb F*�l�S�̘�z����""��	5��5Y��㣣�A������b�]{��9Z|5��=-}&����a������@]����=��M�lt�����{o"������	�+�X�#1Wj�^��KH�P��}���>?!�7�	���f�Ny%Q>F��\@P5{�0?�����ڥ�@�4�d��Y���52�����Zn�;t�7��q�ӯt����x�+��x��kBR�bO�r��p�m��&�j���V���&6��3�,�~��p�OE���@'6�d������˶����έ3zz0�yi99��j�a�\���V�r'2@BR�\&��s?SSS'W׾�9����1����a��
h���)t҅��x{��i�P�؀faW>�^E���[��3��0���;�)�8�o�~7�O��о �|
�����x�l���,g�����P�|�i� �i�u�wR�X�A���!�D������Uν!�G[94_np�@ y�|���0�\5�����Xh���D�܃�uW
]U�߾e�͑�Fp��N���k>O(�y�~-(��ƹ��q���c��i:��#����&�sE~�Ĉz"oP�S��q�Z`m�ͱ�����������"� X.,��Դ`.����j8��Z%.���^�����m�,��\R��X�؝�B������NV���͝O�$U޳�����4��W�83��_ۊ܎�<����ӽ1�#'ǑJ2>Z��<�-����|j��<jG��ER1~C���ڔ�m�Z��>ɂ�[�pQv�1�e�D���Y'W�N��&�_�rq��]Q��u���O?�?�a��/�rlt��
�0��k��z�+Es��
���!JI�A�	���c��qrjj3���n<�@/�==8H_)��&�p�&�V�&��r�������F�
��k�v
�pB��T� �� ӊ��VYxdhp0Yr#������4�����]a�����
LqIIߋ���ѯ��uzKAΜV�j��
�I�����w��9M�
S�$S�,��_1�t.S'������T�֐�^�z������	����������+�[ih��Պ0��j6��2����D��!PM�����g��YS���EXZ�������'�5����gh�,�{�|Ҁ�xW�^��4孤����D_٬�Ԣ{�n
��^zNkZ�ƫf�/RBqY��/�/c�h��z��v�tW�������Q���WRZZ��V�0�ox�����E�֪�a��^�����\Ta�V�G>��Ê��YDݶ�7�U�f����..�箮
���7��j�s��k�z����, w5KNV��4a�l���蓶�'4�1oŻ>T����� ����Q_..Z��?R��{�SsϋSs����TيV�����'�@`��rd��D�\�����S�V�+���2s9U��x��(�����F鹽n/�A��!:FfZ6��s��q�g/*�a��������;(������H�ڔ��F*)5�х&�E{���ZYZ�#�g�_e}���Њ��R�����&{��\F%��z��J9��ck\||}:^@D%F��p��[Ѐ���Hs�����Q��n�ȣ��ô�5���q>���[)�R�#u+/e�q��Dt�>v�Xz���F�}	n���hɴi#,��Ʋy9��C���?�ySW�7�57���1����3�� �<	Xk6���hA0ƇE��DZ��3�0#O� ~Q�8=�_�bt�>�v�ADMM��+Ǟ�[K?�۵���UD� ��9H�k�W}����(���Y�ؠ�����	Y��~z�Y��\�*��"���jԡL#@�;��G�'uΣ�3�S���U������L,,^���a�J��� �����<~|��TS���VF�ݘo�G�ƚ�z���jߣ�	��M`��Z���DJ;��S���+(�U���ߚ9��My#u 1�G���))��UTT���t�X���}��_E��x> �<f�͇of��[���ײ�Fge[| vD$F�'������R��hv�De �u�x�j���j�j�:�boP�.ij��ϴv�B�E�)S�����{L��b?��x�GM+Ԃн�V"�੹{+A�����"�9�Xi�W~�������Z���9e��2@"@�9=��B��$2�}�qYÔǣ�.���yV:�ޟx(�d�.
�nM���(ef�Bh����.,�|�g�ں&��#cK���bqu�V�N��\��gqql 2�@'��[J�u�HN..��<<�I�}��Y���U\�F{�K��[��w�T�܃�s��l]I2O�W$D ������τ�Xmd���ˏX�v�M6t)%WD��]�:���� �ޗ��D�J�5�#w��ź�{�j�S���.�ړ���*�&�u,,F����"y��M|�N�`P���8�a��jPq����-(r�Z���Ļ��TaC##��{�]X�|}�0��;ø��� �<���[*�����<�0%��P���:�S��^�;_��������ȲT�Do����V�ogUz�A[RRn��!�hx4�Q�N�β�Zh]��| �X8��C�moz�{���h����k����������#�éiy'33󟫤�H�4U0��޶���P�|�}Krs�,�M��-��T|�b�U�	��B��.֞��Q�!�l���1���T���eJ�v�>��KL��W?�KH8:9�k��dikk@E��%`<�^�-o��@7T���m����έ~N�C�zQ�X��}�N�Z^����8&&�`��u���p%u��ř�}Ch��2[����o�JJ�'�^���7�#����>y�(��U]���X����1���j+xOD�+@��G!C:�����񹦔���"�NN>�W&$q�W�W'�:;���"��9;��Ղ�=��گ8<�Ijp����N��qJ���H��&$o*4�0Etq1���&A��W�ׂ�N���2�N��漇��_W��U�9Sz�ӧ�~.���ލAl_NE��s!3��R�>��|LaQ!g���HХ}�P7�A���`���1KP�\ �����,�j|־�m_�";����C&�0�����}����T´,"������^7.xF#A@m�@����G2%��
��˯�٨�h���=+�W��x �����%���(y�`UxI�E�[�����h�k�R5XYYY\P̮W��������� l��,�~5�{�_��Ƞ��_�ȠJW����x���]��ߙ�lӥ�k5�,!��Ԥw�j��1-fqU-{;����7�o��,R��ŋ��mT�,�f�Wh�M'V5S������\���MRG��95MGP��*�J�-\��ÁޖII��3�{w�Q�oջ�B)��"-99�6��%PC�b�r�2I�@
��|�@s&�G�/���1O�}!uT��(;��jPD`~��[M��g8�u)��?E�X���yg����y�Pٽ�v����A�T�:b}&���A{mmm�Y�i:�����pXk[G����H���`��� g.���[7�yy������gZ///�e=1�T����|���=�K:���mР�Q0����{�5��.+M��-&�@Rw�݉�)�ʄ���w3�d�DvRO5p���th���Uh�d��xys4��M��\>�f��?<\�]��Y�k�P���i��!�����|�}H��S�x�%��_�~y�M0���Ϯx�zp�8�M�7o�� ��L@?�x`�ϠEx N4�I`|��bȫ :%*E�M=�a��Ӷ
'-�dz����@�H?�����Ĭ�]4@�����V�A{��b|Б�jAw���;io0��x��ҷʩ}��ā��I���=-������;+ |ՙp,B����'Yގ� ���hwu�Q+´P�=�����{rRc�C�j�j+M�X�����T�k]`}>DJ�r
Qo�� 4�?O�'�խ9㶴����n�o@��^s�j{�rek�3�*���eJL�@�=ff153K�f�__��d[��1g���ރ��hW<�,��e��0(��^��_�RR��2��bb���������i��^l�XR�0�ｮv�rY�W
���	����xjb�E�����DJs���vM��S�KG`��h�/�5\Qv�j��UQ�s�W/�&s����$��׵h��ۖ1��j-#ݮ�Cn;n���xA�,?>|�I�~Q��q�$B.Rq�|��~���k({�^i|���)dė����h� ��C}�u�dŚ1��fbfZ�=3��~EC`�����P�3��D{H7Qǲ��u�Г�.��Bh��zj��h�o02�4O�3��pGgg��Ӑ�.Ӡ>�sc
`�.����h��ϾރBͯ<�)���A�*��9�'k�<�rm�:�DҀ�q�ݑ�t�pv(+-��r�$m˝<��m�=�{cN�(�f�/��@��wH`�W)�KI���+p}E�Q���r�j�R=�ԤfL]fpF��ݏ��0�_���ms �4���������1V�z��k~�qm��`�Y[g��R���r�t�E5`���K�9,D��*���n5֌ޤ�`ٝ�u�Α Y�=85�3]\]�%�e�����V谬�tE_�kKkk=�\UF��%@b�44hQ�["��Q�����ktx�#]��D��J%������ft���)'u5��+�|�WRRb��w��k���`W���I�fcph~-�����������MM���"�����&���
9���Pq�E-� vܻ@�}�zj������l�+� 3͝+��;)ꚺ���U ��*��C�
�|�d����B����~CqH�mi0�U^__:S?�+P�c#����s@� X(F��>�_O���$�}T������}/������@ې���lK+��#�5�e���)���^`	+�P��>�ޛ��
�S��\̲��Lo���T��iq��)�� ����X��6���"7�a��,��b�R��?�Z�:|ʹ�e��;)Ė;�ַ͑bc#h�|&�|}}��|��¯�b�\b�/Ў9��EL��צl(�ͣꗁҚ�a��B�7�aU���@ �$�/t�4��K:��m�pv�1���0f.5+�]����w��?�{�PTLl�qD��d��� ~.��:��,m��&?]�P�+t*���ҫ���-qҥ������r(�fߪ�x���_�~��9�Ƒ�h��>>���0>�����i���]Ɯ��ۡ{�������LR
����t��JGlV��#v��*������X@;(c�;вK�2��MǬ�5�Tr�07d����.zP����"eTY	���r$��(ϥ���={�U���>0
��C�/6�QaO?8�[�#�I7j��{U,-ο�V�_{.�lLfu�L�q��ʺ�]D�a�[q]������z�t�������au���e�t��+��jVaTM�"�N;��* �5�@���m���� ����I�WB1Z����|cj�)f�i7DN^�\f������+������冄\5�n�n=���I� ܞ���CQ��R��|�	�$G�s��0q�4��L#��qqq�++�^����ј�*���VS���F������gttל��D`�۽H\����N���H�==�C�%$$�Ӳ�l���N�.E"��|�{���.Ćª�o�;Xc���7&�6li���Ӕz@髀#�vpo(r�>�174�p�2��)j83�tt�4�T&<bH�\UY��`�x��@s�_�ퟙ����q�l� *��ފ�����MQa��Q���8�q5K �P�,��\�s�1����;>�q�/��m\��4�W ihh�'W��w���Ѷdic���������]���oK}��˺
�p�%���H�����+ `�ެr����**� ��/�QӃ��*#�1��5+ P��^c��Xh�Z��V(��߾� 겖^�g�_GT,���|}z�fhS��"�ଘƱGޛ�����t�ɋ�PYi��i]墼��|�b�x�2�<=+Km�4r��D$S��8űwZ]��-�����(�!^C��Յ��r�c�[x�j�C17�]�1䴗��m�/ի� b*���O�u�lG�5v'�9�y�����d�rs�?��t�>�Ӳ��oSX5?b���4���Ǐ�6�~���tn/�5k�;1RNkc"v��fKϝ��ȶ٪7K�,=}d�����W��`����^tIq�m[��>>^���b�X7��m5�R�!�yx�������f!;Z;��SWA*���w��/���ŃSX���͎�>~77��70	��x����B�\��7Z�&B����=��J��aT� TTwU�"��D:�T�U�"�UJ@QpE�ҥ)R#-HJ�H�  RB� B������=�9����3�<ϧ�̝��9���V����i
z� rO�X�~f~���p����w�;���acN�I�������l���ٻ��<��H��cd�����o�ÌM}�����]M��h�۷����X,/\�|c�������>�uwF�7nN/-���I��>@K�ֺ�G��`^�20X�? ���<q����o��"��{/��P֍�:�D�,>����j[X�>}�I0	{`e��|����ۡ�*$IX�ms����ݾ�h�����(erwsb��q���%�m���ħ[�:���6��Hľ�H�������$ܗ���&�]QV��ؑ��V�P*p��w��k�r0�ި�?�w��Ӹ7ο��k�-��4�R�5��:��؃��	Q�����V�N�T��U{ͬ��/���#0^c^f�O��~Ak��uy���a����7e�ȯ����XH7a.J�pG�#g\ϐ��(�����6�����O9:;�J�Wp�5iNO�(ݛ,P"�<Q�����[�%<:.��Y~~����m111	��b^~���y�zx���t�&������X��<Y�7��mT]z�a.*Woz�!����:��`�G)��2O����w9�o��t�J9[�]$v������T�ؕ
����(���`T�|��� ��,z�dR��Vu[\�����n�~���Bi�Ww۴��cR�����DcӀ d��%�O-T"���iP#=h��X�G(Ƚ�p*�4ePZDMi
�ˌi�a$��|���9������X"�%�H��I}3��(�]4>nc�u�gfF�>}  (��O�@)�W���OTA[�eWKJ���
�l��1H��_�!lRâfm�ߤ�پPߑ�6WW�Qw=ټ{~^_]C�� [3�y��֖d��o�"��ȧ��	9<|(E5#��Ln،c�$ew�K�:�,{&t�"��Ǜ6S%��4Zk�fY&�W��x�ӡR��!s��Z��hm$5�$n��A�l]���r��3)p
��|���c��7��u��G,�P5�y�8�Y.�����
�<�b��
@{��| ���+G��}���h� E�
W!k1;`�|�w ;���b���O����_�Ii�Fӗf ����h�������Z��%���[�.��嵬����gT���q^cMː��.$��.�k�v�NN�˂��y��<�j!���y�SJ﫨�
Wr�HL���/�n��M���C�E-yy��Z�4��9�/��'!I�J���r7���\!��V��ޮڊ�YX`K;��@��AN�S�r_/����?�1i�!�9ﷷ/�~T�C??U�F�W}T��VE��Ң�`��Hr���JuH^�{�7�[ec4=K%ư!y���!8{{{��R�;��O�[�c��@.)Oe���{^��fL�I�a��U�&#Eރv3@�h�!0��ɹ��|j���gf"m~[�(�u��S	�9'�h��\d�7T��-�}MH�P]٥�� HBS��d���߂��Fv��?:
�.��rf�K}_.����ގ��xy{;�;Rf�q]�,.�/LT�v@���&�2oqѩ_�{�DE�-|�4楮�jR��h���P�{[w�����I#���Q�*��J��ȍo�7�DiS|���EA�~ve565U�!�1�]V��f����~��2{�Fä,��{<����>B�g��W���v� ��mַE�- ���E�JYȺ �e7����T�.�Tٿ�76.n��#и�mN�!�W럤l��g�y�\Kk��H��|K��wS��2��<�>%.��U����t��p~���J ��յ����70Kg.��ދ4��"0"4��T*�[ӂ��5���0�P��+�R0~s�g˪���8�8��fU�V�p@�.|jM=Y��)N#E*kb"6S�C(ܳ2;w����s��@Y�Cc{����0���HaLt�k�����ꩧ�,HaA� X��_ė���\�IX#��"31��_J��Y�5L.xK�,n7�(��a�\ʮ����0K�������"Wr�Z�����{fU��l��w����D �r��Sp9�����m��V��!^��9�l����OI���4�5��˦���P�����&���d�����_�Z����<G7/TyR����Y�U�ۜ���We��4��(�a������Ll���"�fUQ�E����Ռ#�f�c���w� 1jd��~?(��I�HR��݈��Z��]|P;�kə�.@�I�:��WĀ8ڻ�/��37�N�2#�ڿ����b��$�nD.w,��6�J��;���#s������gf^����{a�
��G]�>�F��X��������}-G2�ʓ叛
~e�� ��#������e!ڴ��I�IL�QBOV뙘�|e/���	�/�jjX�;�qyV���ׯ��)���׼�~���wrh����B3��I�^BCG���19���LP�7'Bڎ��Z0T7W����>C�Z�쵢�N�L�7YG��:��\*9�^ZT�Owe_�4�3`�u������J�d2�Ex�J�T;dw��i.|`�@�����޿ln���d�.uW���t�?R�,,6Nݖ�!�$0��	��d��4f�
���{��-t�*P3V��>��/T��ۛ8�\�pe-��w�F]]�K��K�.9>|hz��u %#�U*���цz�K�
�z��c�ӄ������u,�N1�2����>H3�oG��8��e
MM0h�]�2��������(>�� CL���Ư9n�ŢS�UO��N^ɪ����^����s@��}H�ԗ��KE��{�B�Z詳bs�2���%ҋ�b��3�����\���}��B<��_׍��Ō�g~j��@���&w�hС���(�8�w��w��5L����6ȳtIj�� >>>�����P���paaa^z�v�'�� �)G[?��u"�<��T�H�e`��8�Pݮ?�H��6g��NǢ4c�����2�*Ȟ�۫o���"R�.J�~�%xwh�hHp=H�4N���ʳ����+��W�0v����{��*pL��ϗC�U�2=m�7�嬾��!�K<D�2�韮�
�{�x�H"P�ԥx����(����5�ӡ�ɀ(�@��XX���b��?#6/EC�'����L�&���E02m�����QZ��A&�s��Z�72Ҷ��2%�Kv�tt���SL{=�d%�o��Y��1�{�Ҕ�r�1W�b�k`Z��j� @%-}�H|�ߥx|�u ����������]����������L�A��W��RY�������/�G����,,�.�4�l�6��:��;�7�2���^�]
Hg�?`��m��I��z���bm!n[Ǉ6�"1v��_���#o_�Jn���/��I���՘)�BⰞ+ҩ�>y]���[�
��7>ߘ�n�e7�;b �ꔟ���a��h��I�I���F0ɳI�3�Tt��퟽ v�ֱ@�s����%�����>��v�j��N\�A�$�� G��](?e}��wg�%jcw�3�	'u{���N���@���+��6Y��^��X��ep/��X�Ԫ�E�x�O��V�M��SP14�50ԩ�<">����<{���dE]���}9����-�����`�8ϦDP�I7'���g�0��t#7~́�r��_���P�M	�V 	�ChRQ�7����?�*�I��S�d��쒰
o�U�oF� ջ<Q����uK��(�'�	��4��2Z�ڗV�)�v�Qԅ�������iC���[�f����e`e�-�c���;m�{�[���*	���������)U8DZʰ*�sH�D_9�g�跽~�k~�/�o{���4�/����y��-AYB;qnſ:!њ��q�&�]�c.�h�$�̼�rX�&#mCp�=x��?V5Gmz{/��}~~�Q��������8��X�� 5hc5�������
>7K"&y�6�����n�U��n����Rxe�1�����Ǒc��"���������|�q�x������b��(+ ͫ�a��566u�8���w%Y���7W���q��3�$��>��X{	pߕ����or���,��éd�.�����=0y���&���76�f��-&W'__#]ݨ���R=5TR��d�l���I�����jX1r~�(3%���b��9�,� ���"��Y����n�Z�_�}�N��f��tH��MOgꪶLʮ���*g�a�e�=���}�$P��B@	w�����#�� 	M���<+��/b��CջE�$%F@����CV|{p���ԭ?W� �kt��Z!�`��;x/˿&�R�x�k9������7<g~6:S�O�5h>�vFD�������y/cY�N��0γw[D���_q�:�kCZ���TwS�*�R�d��o[�ޱ(c�j=
��j�2�^<*�hJ�u����1��mm��5�p��H@��6�4[�����a����5���"��G!�Ɲ���6��2�*�
��?��*������o}���iM��%?�x��6�^�V����)�H+�{q�.�v�:�C�����~	�����^���x�UV5+���}:\�:T�9IF�����l�d��|~D��:4�r�ad;�腽`�q��~�(����P])��Ex�=�V��(v�5�~��	�,��f�*_�l�u�L�P�O��@O�� �D�E�t��	�$h?��x�Ω쾤QE�	�������R a\'S&)!g���R.ƒ��ln� b[��i��'��C.���i1�������&��k�W7NPF�
���z�
�TV�Ju9e�w�T��L�#g���ي� �Og��ȭ+�`�'ɏ̀����1�<S�|(~}C�d�~�~bN(��oM_?|�]h���dޱ����tV��x��(�=�_��0(���Ac�j�dJ�7d��]hi�!D��Oٝ'��u~����/g��ů0:�v�*�����"��
E6��;B���v���?*��QwX��)���b+^k����5�w�>�&ppk��_�J�d�*9W�%kP�w�9�?)�A�����b4r&�`�r�����h�!�t.�~[ZUQ
z�N9nv�g�����Y�$"��w�,S����s�$���@��w,��׫��)�2,I+~���(K�*��'���5%N�r	����AN,���.��_9#�j�;�v�bh�xJq�ᆠ����L �z =�c��E�T"H�k@(Xrl��}���O��Y��Ā�4{ '".
t.Mu�#�ʋnkk�1A�ÍJ�s���YC"Q(�ԝA�ӡ<���X���d2f���	Q9�#P�����D��qȳ%GM�����Kx�Q����7WO5�C���$J��mx8+�����w��!y�o�T�n0��6<-r�Z���~y7�� T8$+K�6�+����93�N��T��Z+�:b��F��mϛί�x��5����|����ו��?ip�wg?wx��c+y��ƽ�W��z�t�]��O���
3��Yf����_n��*�b[)�����"�E�U�;�"�D��5�������ɴ}3�0�7�s�����k��]�	�X��Ώq;��7(|J�6F�"��y��dd;��#k�'p�n��M��w��+Y���)ځ���;�4j����#�].���/݄�$U	U��3�,z�vic8�E��_��*��A��&e�Y7) C�x����}�z���sٞ�����bblj�~��"�[��g���o�-��YYY�R�(��`�	��/_�(݉���5
o�cƜ
�v1V{8e����3�y��������ó�����
��%����O��-/��-��$bN��t�� 
�t��s��D]B�Ѝs2h	����U�>yBN��� ��Bq��)�t����"��qBC�hu�iu�Nn�'|�S��F��=>������l���
Z��HJJ�(Q���~��+��[�q���3���V`8ۄY�\�S���&���A��}�h%Z��l���'�>}�7�$�2�n��1�h+2��%N�4*]=?�������:���w�(U#gy0����sH/Ѳ�omC����	�.m�3n�պ{*.(��n"���=��Z�~@�1�peQ㳍��F�U��t��9�,9��SA
t�8ŗ��##i�I���aFg�F��L{�������Uj1�"��ǳK�=4]fs~�֯!v��P�F��6��;W(���v�Ͻ�jЄ�0��s���,%p¨7���>ʱ<ϰȬwaA�O_:��|��F������5�vJ��5e����]5�Ϗ���5���J������v�����m�N	�0����G��GiiU��iߔ�?�/S���Z����ro{�r���me(:����;�Z9���Ռ����蝜��;;�pG�GF�$f�҂v��<h���!������E��[������(«a/ �CB%��f� ����ac���Τ@�C���(Ƨ����� M�W-���_��^P�L��X�����Ӯ4�حO��9BEo���d���������?�X����A�BCò�ڡ�Kk�����}��l0�QD;E������x�L����־}���3/3�i5����m������!�
��+��SN��5.�gy�y��q���X���-�(����G:M�[�h�/�3h�#[�:
t"��Z5?��x2�Y���ꤢ�{���Kp�yu,nWd�B�8-��C�٪x�;�M��#	�.b���5r�%z����;�lyiiԟ$`jyǷ!F�9i��&yr@�t��g�R�N���Omй�b/�Ϡ�R��"�.,z-N���U�O8	�V �a�©^�
�>�ڍ��>(�V��%;�75@5g������!0�U~�61���8��u?�lw��.ޔ��`��h��di�
�63��1X/.6��{�� u���w/}�7�<���k�����S����*iG#���A��T�=y��јV�ڍ�>b_$f�@ّ�����h����C}>��^Y"Yf�wx�B��t���\�<@NwS7<jW���S�7�J�	b�%�k��p�IpÉvНsR:��3M͎)�]J�M?�h��\k��e6G�?C����a]$�k�US����M��4�ڗ�l�M5�h���V��N�T�]kx]�Q���4��*c
�g��|<c �k�����W�J�/���/o�T�u�(��Ү,���kV�St����k��f���Z��R���#ʳ��(v�?5�\�c�X|F��z���������݇��>�on�*<�"�Ku�[����I��7t��=�[lfgf�p����p&�Z�mOƲ��T��6��1�h,8�^>��	�Ң0�i��}MG�I������̨z�$A�`�U�(P}���y�q� uH����  c�IA��M��7w�ړ�1/�v�C'g;���F�7H8 Τ�I��Ih�����VaC���-u�l_��ٝٗ�W����
�|�ƮP�j����1Lx�Һ(|Л;�I�%��k����;���}�k�j��T�ڍ8��br ��4r4}SVm����XY�3���9�P���u��^���c�tU�Ӈ�]��b9�}��V���6��ڰ��07Zҿ��T��_#�p�����>4^.n����u�w�A�"\Uov�.��h���0��>������6���@3���F��b>�(���9����-�k1�Ԫ�R�fT�eI~.�C{}����3�+5C{7g�����@����o5���0c���KM�[	ƨn�M��!�~��5Ԕ�Mh�:�<��{�M�ܐ]��k\�¯�t���ѪhoN�"z?�w�N�����T&�/^�#j�WK��j� �a��-��nf����;Q�g�9z
��n�Ãs�K݋����l2Ko.���A��z�U�)ܿ���f���*�s�Cae��L��q�^�O		���y����:��D�����|~��L+��f���@A�y�����hj�N1ڗ�X;OiX��1!g�؏T-,\�i�|�2x�S��i�6����]�:a������?5���כ�� ��!��Z~(��U���,�X�`�@�.;�w�PrR��8�k�u����o�}�
�d�P�N��X�-���f^��%�7�r���Z�¹�����C'�$C%�n��+T�Y�n� :� a3��WU�H�A4��K@Ԩ֜x�Xd�B�d��C�⟩�������m���ac,9�����m¸���-*h��^A&Ī-��fͣ����J
�,
�5��{�Q�cZ����Z�:�Oz��q����}�
�������|�WF��;TGք��m�q���FI�KS�!G[l�R����ׅ,�tn�s�ʊ�Ļ��6���)mMM���ߍ��K�ؙ�4��眓=��V��md$�ǩt�QK��?�E��2]|)�������5)��q�t�p�C­��ԡ�
��s7Z�+lH.}۩�m䏿������30(4���r���:�. %G�ם��%]�{d ���h��^�`R�TKS�5�#�9p�7�T�ϸ�IJ��!�������?'aD�h^���}*���Q(��N�*W�O�Ҷў፻�Ka�����+4��
 �ne�CG��#����� C<\5�ۏY}D
$�Xsϰ���;���T'ϑ`9,�O�TܕP��8լ:���%�E��eg��}�ϪR��Se�7�;��UIb�kk7��&��ԉ�<��U�b��z;x���N�R�3���=���L4<��K�8ǟ� MA����c��|į���ҋ3%�@ �C"��(�
F��?��6_^Y��b]i�����ƫz���^���
��>�Ԋ#TT���W���\=բD�k1�����o���g'����s�H���N)F�Ȓ���:F
(�Ui�\��]%V59���
 
I��k�+hgG,�h��M���-j�Ū^�ؠ]$|�4��{�C�tzow7H��-������	`R�:Hױ�5Uy�	��	?���B�Z�o�5��K$�_oȱ12���eQ*F���L��`�~n������й��m%c��2�nC�1s9����:@T�����s?o�bB�������{�Z��=D��@�-sFÆ���J�Hm����]�Y>D7��Q�t��d�#]��My�E)��m{�݃���s��I�V�/��Z�0�E۪l�4��?�"zv�4Ԯ�L�ܺ)�a�p �<���F�w�Sn�n����e l�wN�vPP���J��źK���&T�8�gh��C��iW�NL=���h^On��O���-��~�Q���o���j#�DX.+g���o��ɗ0���2|i{���N �!����|h:/~=�C'�`U/�U�]7�7.d��Q_`�Vگ��E��/��|�n|m�9�	�n5�FR�Q���Jm ������-+�q�Xk�J�m�#� ~j����HdHش��b"@�
'��YT=9p�\2U������yhv
��і�YXԕ��_ �z�]}ȧ�W�f8B��f�?�� ��� Mjkk������Y��}y���7�î`* bX�h�Q�$u�n���Cu�!���V�!I|(���V���{����J�$�s�x���8z@|m]]�ΰ(�fC�%t�z��z��/�޼�]�� �\�\�,]�6\��Qw�gp�?j�d��9Eg�>��YMؗ7�.��%ݱX�\��XT�%��(�/`��(wfkk�40G�9B��?�C��2�X~�\���*Ԓ/��}�]��v�a��U.�mmvG�0c�ڙ�Â-��V�<H���6aw��G�ڝǗ��.�w*�%6[{�m��"?��Gfe)��.�R8�$gx?G���|;?%e8��PT�Y[/f$%��8��޿G��Kw�F3��|������E�����PM���O�t�2H�˯]s��#1���J��P}/`PWk$(�v�G浵������j�Hf�# <�fgmo� #=���M�����\u�查���3,TF������zJ'�fV�4	d��Ɔ��?G(t*�7�n�vt*��	D��/��+<�_�{qNyr����b�1��*�Q_�[�@ɝb�c�������P#D�^�d�404O� ĴI��*~�r,��t�*v��#!G'����
�=L��mI+��g-��K�c�� ��H8Vh������Pҕ�RC�LP��fP1�%?Z�kn�~���ՅS͊� #�X�ud�(k�����[�98�,ȅ]�% u¾���� e����v��: �&��JpK$����|W<3�h%ῒ�Lp��48X`�;����	�(���a��Ԥ���hլSmN����.�h�j�Tr!06F u���<��<	͋R�_��LL�:�g@Ӣ.�Hzx�^�v)7fأc����� 7�<����|�`|i� ��̴�Ք�@��������&���;����x\�i-T,��yؙd��=p�(�^2Y��u�U7___��U^��Uk�)pZ�#�fY�ޝ|����NF}tK�a�ן�i���-���d�P U���q��������kE��

��N�pg��o�7|��N��ƕ�L�bE����D"�ɓ=w����𹅅�x��e�6F��-�>\)b|�#�#k�Q�<GhT����t�Fj�b�'�-����w��Z�?P��Bh������;��&z���+�w�Z观**^��#;��/�ɱsm�7ط�hyi�ʛ����18����
d��1�Ċ]�����)�ij�AG�>n�h��!^����s!�i�U��������M&���G6 t����g+޲q�e �R��3�kg*N3�-����9�k��������_CB7 '&^ �6����@-��T9Bٔ�lV�{<��\*����HW�]����`�t���l_��iP�ڰ=��"%U`ꢌCV,o
��՚\/u�} ���I�`"*�$T�vl�B�D����Y��#�k�}���~2����6��1��w��֏�uww������#}��q�=�ov�����m�-Kcg}����J+9e�����r�L�bT���L�����;{��uw�����n����UV~�z�Ư�=�[l��8���X�x��M�M��=��mq���ӿjg� ��@L{�/(��#B����ʽ:E�z܅hc�ĝ>@e&&���~4ٵ��	�lw��F�־B�	���tgE:����p�h۬޵e�rc3e���v�`�j�����2�<:���>���9��d���#!��Jl��&�����t�������`�3������o9��iQ�	j9��1�'�1�����"z�y�4���_Q�����{ĳ�~#�jo}Kh:�3���2677�l�� P�֐H�����qS���?���ݟ�����&��QW�~B�;�{��P7-�mycr!��71OJ�0[�u��N+����֤����`}>��O�V+K ��ȱ:>^I	�jR��t�n��r�s>�ʍoL�e�zI�^�#�䤧���3�_Ct�?}d?�@�,~N��Yh.5�1�����o�� ��wyܻ[tyI���v�0�!��-*��e�(�}���|��б��k(6�B��p�!�5���s\�gz<��h\�lܰ�j}ܗ�t<��5�#?��XcSA�a.v�:ᐲ�������:�&�ݝ+܆���������כ'h�r�B��1����hAD�	�͢��)g"¾�@:;�{x�w�̚��4o������`o���lj�[����8���Y�]y���%)h6�m6�a&��z�f7n����Y��ڞ#�%^3F�5�.��뚘�M�VJ��|�N����x�<'g�e�
�ڸ0������heuϒ�z��3c@+A����lB1��b�e�Z]s�rNs�c�������:m1cI���+��;!I}񥓢�oc�?އV_�g���1�sQfg{�����k��J1��x�X�����cSZ|�İϕ�[ǭ
��́��c��+� �[��Eu�,~������T�<��C�H��@��I�vk%���G聃���'+&�f���oj
���]�4@a����i��Ax���˖j�j������LLLjV�A�����S<���|Vw��l�b�luzp���ѣ��g)�;��K&��S�n;f�)����Ɣ��WIM�2��c�N�K!eP'$@�6v��`獵���P������#t��C��n9��>8%/�Đ��P��e}(��y��cX��뾱��}�,��Mw�ւ�U�jkE������C5��V��ho@? ��ɩfc{r�bF�c������?�RA%zhӔw��Z�M2Pu�p\`)ewWd����S�X���P-��]w g� �zM��ɃL��UT��ͤ�ٚxchtP~�66F��&3ǘ�Vm'��X��la >���8s_���q��ͅ�����Z@.Z�(ѱ�����o��ola�[k��|JLT4�~h��-�ҫ�=T�B,�9�g"ى�e�&��2f;�L`Mdl�����L+�����ݟ��+*�RN�^ˀ��d�������ag���@��@ޑ���P�
�v������$�#��tFWo�wWP�@gy��*�vTy�C��.�c4<3���ʹ�vsҁ�^�xʉT1Ћ|�ľ�؟��#"�����[D�i������=�z�����g;���H�ӷ�|�b�����+��h���1�X�ʼ�Dq�]���Ȥ?μߧ��k�	�C��&����o�Vy󹊖���!%v�����[*�U�*�P;�a S��h�Ym���w2#�����<>����w�	����$m��?�i{���E�����t$8��%y��Ob��\ll�O	N�j�.[�ݲU1%���/h�s��'r�T'�����D�]��<�>k�'?�~���꺕���Onu�&*f��$���a�?�ح[ �%�� )/))X^����Y%J}�mT���:����g��/�`p�1����)�W!*���u��CY*�c��rZ??&���8B#GLj����83t�TKKIؗ�ݫ Y-l�PIJ���!�n�UYD��8������Ą����i�}��y���0�諮�v-�Y�c����{Z�Z� T�DG1�6��O��?$�^Ze�O��k�[
�$�+$1M!v
� .A���DW�C%P 	�pHV6hqߴҴ�B�u��Y��l�8zG'73&Ʀ���ZF?E�¨UlD�rMX�r��I>��n���.��㛾c_8��=幒��fy#���])�I���T�0$������5˞�ȍ.���Š:��>p�b	D@O���H7�>�t�N0��L߳����^���u�� �cwT��G�����e��m��e}%�ɲA����09�,��o(�di��C<�ַ�s�v��=�?=\n�~�z+�~����0�G������\��\" �'m��r��@l��^
z�7�3�}�< �=d���`�,&�Ͽ�ȁ�A�qB�g>i��?�9X�{����sGGO@�k�]:։����C���CK���c&b:^7��x��B�҃�>��*�j>�%��,��ω�zh=|��`|�CB�?ڢ��w[K<W}���+.�����͌3��������ҟ�7�-�'�I��>"�=Բ{<���Pg+�1�ogGDh�S\�)9,ջ�ig{�F�
�H�h�]v�U�FA���^�<�Ψ��A�wY�����Do�@�Q������=eD����T���\�n�bB�8�����3����#q_�"@VfeA7O�}�TW���5�_l7�aqj������錇���Bem���jKLk�{6&%-`�xxx�-)Ȟ5�Af��_տ�=Z�&�{t�k|�g�=�����R�^��MF�bu��vЀ�1���ɴ�D��q���Q��Ҏ��=K����67=�Zhs �.���s'}���KG�![u�>Q��]��-���G���$H�+)x�(���f�(��)���Rn�w�)�1$���k�I�մ+\��:�>}J=�u���;n����f�� �k ��x�e� }��h�N��A"�y � ���1lw��Yj��u8���hC ��O	�i�ӵQ��&'��o7��nL�% ��rs����n#ɪYPPD��A}��� �N�:�b헀s�4���3Jw(!A�սE�\��?`��x������nx��72};���w�I���c������x5�S��޾�F���E����t���
3`zQ�����o-I(��8`lf���P�2���	��q������i����C�Y8.���Wo����s��_�2�Z���3`�<��������n�ޅz-���}]]��� �{�i���F[�@?�R��7'4Z�)���?G���g��=�ˁ'v� IA'�?a�JV"�.��c��p;������H���L�c�ss���x�Ԉ�x(������!9Lp�;�ZRR���Ϝ����s�I��f�5���{���ai�xp�i�����WJ1!��������������%�<#���AA�v�m��"�.{ػ�j�=��BE�:F�]H�����?���0�P���[d���N~���M�[������U���A?�1�$?���^�X�&A:��(Vk��0E74��'ï��.*#�����;�U�n� �j��"I��9ձ����k0ļ�&�И������)�˿tsl8�����TyR2��q1��S��y3��9�������dp��=x�\������}���#07	xE�6#����$�r�S:{��j�����;�K���P�9�1c��Ǚw.a��ۿ%u�t�(U�>���Aii���+� �UBJJ�����߱Q4:H���?��@�����IHJ�����3}���&Tp����Pu�9���7-e��h��1�}Dp/��N��"%&Vh�*y�[����ڻמcM^bLi�,��_���α��{Ȱ�#��$ov��IIe���d{;fbr�������'ؒ�xQ7�;�
{m�#���4�՛�����6���Bܵ�H�r0��/���!��vIW^�v�� g@d���e�P���" �A�r����\a�f݁2��3�	�I_@�/�߽���(��wm�����F�	@�D�:B,׀�=x���s%�у��Y��탶�l-��mHf|������j�d/x}fH��:���4�������~^��&˽BB..�~���aB\di<�L
lZݢ�-g�lы�7z��I~�g[��o�y������-�
��@��w�X0��V�^5�%�	��j0�� ��2��{���������������HD�t�޸�,��������ő��ِ��f�9fL"s&��Z[������/C��<���~l�Q�-��,�=(r�_ �媭oI��_w�t��)\D�#''g򂤤d�nw�K�1QI	��!=ՠ��{{>��c�x<�[��[�
�KU�C����/��)�;K�1�
���A\��3�+��� 6+ PMW�{zvVz)��Q���E�:�!�O�� Yq��Q7Ru�	O�&%�h6'I�[^��bKٹjSzpe����IJ�٠��鐤�r���hxxc-�/(�y�lw��B�ԩ|8�A��4�����9{DD���x
ԟ��Q_C�1C���f��15��<���ql�Qٵ'��������������0?>:��۷�P�����[����#� _�:=K'����+��6F}�+a� ��ˍ�: 髞#I4�����]!l(�:p����-�ye;L�_�¦$��f*H9��|���Sa'���δZ�_�)���de�����2eM7��x�U����5�۞��?Ѡ�.V��RKl[�ْVv���,kf��8$����y��_Y��Qʱ"�7�/N�P	�����.��1x�g���i�F=�Z�� mѯ�nzZ�fym���=z8�|&���q9"�k@q��}2����e'����=k�1��ץ͔�o]j��M4燹�1q���������:F���,Zl�wh�����R-�n���F����~v�ш	�X,X���5�z�/B{�Ą��ޣ"����\��K���� �Ꚛ��$�`�([9�]C����RGd� `�}���A�}������a�`D��F��TG�V��4�~�����Q�d	/U4z�� ����vq�u�n_�O�X�a��0&�fA����
`%�
� �A��[;Q.AC*�Kr�ah�q7�"E��=�[K"�����o��ꈲ��z�9�f�O���Z�h�"���'��;xmct�������Fi��޼��T�\22��\�k���n�����D�2Xē��e���i���:�[��-����H��"�چ�Ln�bm>���Q��y>��@�10ЀJݯ����#p��GD�P�L��O_��u�Ի�p�v��F�T
�Yx�M.�/f%k��|����\?�/���pK	�p �-�V&��j7nY\=���\"�Zs
���٪���
����B�eJC�;��0�=:�L20(;�|T���u��l�\W������a�<t�.axd.Ĵӥ�^6�������Y����ڸM�3"� �P��f�Bp�*���\����S���:���	ך�{tp=qp0	�(tƫ�Z�ʼ2<ʺ>��d l� ���%�_QQ�U9/&��vy�Ѭĸ7��{<�T)_��ۗ��S�5e��t\��s�ӌ���oY��d�����?x�Ů�y��S���%�r�Ue��>��p��`�0%O�ɍN	ڎ}ӆ�|ߤč~k�)q���?�R�9C�]�z1����'�׫z�q�l!4������l_"=��3Ր]A]��d1�n|�YVkMsn����I`��:%�mX<��$�J�t�]W��4�U�EwllL�k:�T܋H�6��9V�&۝���)����R���Fkzxx��a ����$�#q��9���@N�1c;�Ph�	�b'�Z�m�w��j�|����d)_�ܞї������pO��8� EM�$��j֚w�4���T
{����W]���~ඪ�o��\�鮚�7�:|��P|i۟v"�KP����mn�WV�7�5䏋�=='�ڵ��L#	�O����f��'��I`�t�*z�N���xn`D��P�7Ѕ#�4����H W�����K�ʪ� {"�{��
�v6}��#�|�e���ۧ㳯v��M[݋�if�ǵ6���p�����8Wk3��<D�#�޶N�k����ШZ�Y�|��3
ڙ�#�,K_m�C�����j�ҁ��̼t���{8�lvV��6�E�K��N������o/��'|��*n�\���>JY兕���dV�H�ka�;R�Ŵr�Zzc;J�J�pb��k5����`�����0��`��)�@_^����EHp"�$�x�Ʀ��v��msɌPL��/���S�8�`-���:���=d��gR
"�;��9�w�������wqP��C L�6���]<���v��I�h<m�JXƾ:?wwU���(�yOqq����2��(L�š@OV��R����n\⻎�]~��OT�q�!U�{�bT�V�(�۩\��;�Ǚ�Ha�l+��)��պ�I9<��2��O�ƞ����UJE�#$e����\���cz��m���,6���~���]t�/Pbh�[���g_ZG̙���uȌϯVYme���*��������g���^��"�B�Ԗ�x\z)�o������c�w�9{۹����ʅ.%Ͷ���ZK�*�o�W5�����M�ޛ���i��Kwy�څ���7�MB���P�%�������6Ck�����a>P¼���_���s
�]hPk�#�=�I�a�d�}�`{I��;�?����o�����h�_���Cx��<Sh��{��<�|����ⳳ���
���t
[ZW���4_��Rv��mv�)�O�e60�2%4:3AUk-�E��e���:��@��كG��[K�	��.^,L��f�n��H>?�L�Uou���O+ZJJIH���R�]��l�g�[�D!�}�"KCI�ck01J�%�c	��6���}�.W\%s��>�����rP��\�]�F1�f1��1���{�*��Q�ϛ���o6@pfB��n��:֬t���9�NGEG�WkYL���kk뤥�
��
�)?�$]���9r�Jd>��FR��-=P\3���e�~zSh�+�h��d��).!Q�������:�yI�{Y�7��`�� ��,�� +|�����u&�!"\�����5�-���_{����q�:����b8�Q[���hx���;�(���F�H�1Xz��9��s�"�����Һ�.�
Hv�������y�����`��#�D�V0h�Z ,�>��5��(K����76A��@���i���b�X�aVȢ%�N����Iw1���t�`��ݫ�,;��̻�[e�IT�� d�F����b��qɍ�K�"���]ŕUU��-KMK<���1Yw�y��y���7+���^�!�t�u�
[#7+�����G[�Ui<�6G������^�5jVἡ� K�T����1-�Õy��0$���/�l�毰C���� �b��������V��W1|mg��^���L��:^��h�/�w���,�|ͯh�N'�Q�ւN�P���=:���q��Z:Y��o���x�g�,|9���]`�������-��
y�=��ME�u�H�m��|mb��������B�K~b+26I<K��4{�ۻO1�uX�J��Ǎz�+y ���$������А@�

�u�v�. ����Vy���.�Vw�?�:+v�������ՒS��8à�\48XW�u��ߟ��$t�z�}�~ e�߿��`�𻤜xc���^��V�k�_��?ج]:ӎ1_��w/��ݲ�^��w��
>?쫝��m�c����/������=d dT2�pG�C2��s7���˗/�I�G"|b�&��G
tX��v����3Ul=�����뽏��Y���G��**��hu˭v�����|�M=R�+ ����g���/ķ�³��HW	@��E����S=�<W=9h�������p����������I�h��1�e�m���F�U*���~:�� |N��^k��0��g���]�
�w��Ƙ��=��r��Aj+s���$�	�_���y?4��6�(��%��C���4��ۚ#�ൔ�7gR�s�V����c�/�2m���󹕿o�����%�����0��36�hE�-�[��`-2,.�oWc��x#�=?r�w�Yk���΍���q��9�.7{�5����h��B��]k�Aa�����*�ߚ�u���*��|�����R6���xB��$��g�B:l�[���%���B	�S	F�z�^6��b_�G6�ȯO[���)�3R�<�����2g �hDF��?T�=v��۹x����ju�T2x4���We�{狅N�Y���q�ji!vb5+N�%�Ea	�X���ג��
;���jp������.��CϢw����^h�k�)0(�	�����x��%K���>T�s<X{��&�sސI'�d��8�/��K�z��Y=��w�}r �$zJcg�I����i��q�y!���:����5��p&��~U�ǫ�˼PMk,��x� @8�z��iJ:�J�w^9z
���Y#�����"�\��y�����h3��Μ�R����|������ʷn�je��
 ���Z�L�d6��Ae�AL4�]rnkٵ@8��`@4ud;�%pU<��Z�p�X8s���Qd�!d>�]���T�P��
r�䨟[z+����~�7k���'ૼi!1��>ۯW7��.e��d���g���y
	���Y;x;��%\Y��&� ghx���v��X��Ǫ���qY��dt!���_�<�,p!W�)  �7v~o�z����c�*��b��= Y��4�ހ*�V�A�tP��3����T/$���(꛴�膺{)a̍���[��F|SC?�'@1<��ϱp-���J�a�'V�\��Yo���y|�Y�����J���i���'�̑� �rtu���I���2���o;Mn�eGG���X�{q��牕=��J-9�e����՟������b/�L�+M���Y 0�����v��7�h��?1�W�B� �ƒ94�}|���ﰘ�!s�3Fv�#�p�E��p�� Iv巏�=\W��3K!$�p
��+{�ĉ����9+��1#2��$[)~��W�졮�Wl�E1��37S�{��l|ۖn!Z���7k�s�S�A���>��{n���ɦ�����f���L��W�ڤ�\\\&��Ft������WQ��J�fZ�9�V0V��)�]��Z3��;}?�tZ~f=jr��f:�-�+�YT\����/�g�U+YWhVS������`;����|�s�}��lVx821�f�#�",��.�/�0^,��ƣ^����;1thb'�%Z+���z�0�;��\U�p�Ω�1�F�?K�{fsss,z*"��W�y���1X��l���g\--���F��xUF�F�cU�����!�?�hQ��R��|�t�!o��諀?�ƾ��bbb�l�0�� �2��ʗ����Ɵ��������(�fWś�#�ֳ�g�;5<%�}��P׈��I�d9����7��=�bo�>Q>�����V��ipAn0�IB���+�K�-�s�vv�]m(Y$�sK�����ҹ��/�S6�ee!�:�������7N�9N��R�����NRk'��S��Y���s>�~��N�WWRr���4nsjȊ� XՏL�țl�B�s�{j�o윥����d`}����G%�x�I��Dֶ�||�����u{"ӿ���,v3ڰ���}��5$��i���������)0�C1��h�^W=�S��s�O�c��>�H���gKi�?���4Zo��kk���e�j���1���lp.�����<�)��6�o��9L�+�B�	^�S���b{�e&����Q8��Y�ɩ��]���|�1^^r����ĉIj,[n������tڜ	��<8i��-&�m���YWW#�:�ܣ��*ccc'O�Y�m�`�I��&���Q�.Kos*�jG �D�Uz�z�����!�{d}v���Xl�7n[n�b��yT��Bl��j�͢򒷗�������]�3hZ�$��o��&�C��R>�=��FaBI���H����J�)�ɘ��>�1���APr�V2���?�k{!d�{��U�ܩ %�C�÷��0��QM'B����uM��1�Y�c㤵*@��ݕN���龆�r� 0^W�?�
[ܤ[��n��RFx�c9�>��r[�
�΋6tQq���9����߾��r�ȗy���	���o���UT�N�����'t+��!�@��f�n��j�2���iii���[0e��d�|�,G� �d�8$2rǛ��~�xc;B�y�!.+�]0N�D�_Ѵ�wRCN�v;aXPW�j�4�]�u�^�}M�/?�Y��<},� �������	�X������|xP|W*炏�:��]ڰ^!ZmX����q�b���Ą�F7ʌ%������
纉�t�C�V:mSĞc�Q��Dے�ox
r����~��/{�Y
`7_�|FBJ�w��=r�]ss��A3�����n��浢�h���wJ%ee��G�N7� ��t�����Ip���wt�]���C�b�r�0h����Β�� D"q�D��Q�t@*:��ܝ��)�~����"�`Y�|΄
��֚Nn�F\޿����T�R�a3R%*�u�oy���->��1~�\���!�P�L�V��k6�'oʰA�OO����N��t
��:�nIR�<0X����kǞ$���dوf�O+�Q���(����Q�\]��DS@m�\]���K�^���%�1ƈ��jv.]	$��D��ՄL�a�R]��ع9�T[��ϒ�)�d'2�{R\q���}Лڒ�f�B�X�����_�=����&:���6iE��@�K �[!`���0J�̱��is���u�q��N�V�$u�uvuu��W���}r:��۹2	�F���.1,F���M���B��@�2� �w&�Z��8�i��������?b�Ɉ�rD�� ��ԝ�v��2�2T��������U��z�L^Ǖ��޸$��舶�>YAV=ooC�����8[c�Z��C#�������+eD�=�5����!5@�N�[�5��V����qa����e��OG'�8{�$ H80`nʞ�YdwGn�w��XB��%)ʼ��%��z�-��Fn,��Lw����"�	[A�~�h�`���O�숱�*.���ؠ���=]
����sso�u�T��!�JK������F��z�P`P�W� ��)�/r�Gi��##C�R�.aH�0�����Z���%�C�
 O�F��@���3��c�>ux��� ��p����³��p]�g���Gk3B?ѵ!�I�^ �x����3T����f%R�L	�D�Ϸ�K_�>x���� �¥$5��աX��F�j�!װ�&u]]B���<3��ܜ���)|,m���$\4ʃsJ7-1���_�82�BE�DP6���"�(�47��B]0U�q�O\��B��n.P��7�.΁�4�n��͝��K&�X��r�.�b;��&5:�FB;���94��V���eP���4?Aۊ� pI֝���pq�����������2
�����ա��dj�ND��']ܶh��y�$�ͩ#Ҏf�܄N.�G,��y�ݛ�t#��E$��Wy��嗣�=�"�(�#}����7��&%����m���b���#W9��ss�E[�{C��8��:�	=a�w�a���,���x�ދC�G"[�k��a�Ļ];t��L՞��,��tG�Q�QMw���4Ҕ:�P�fgV�5`������ǆ�ZhW�R����B����9_������vuyA��ó@>�VihT���! �u򤽝�)`�?c7*��^���#��������Y�=�,�:<��Q���r�;�����#0��	br�*�fo��˲Ȱx�5-�A��3C�}���Xc��4��j$&!?����wᠭ+�Z�:$v�ā_��220�J��F��~ȓ�V�����k ,ȗ���,B�~;4<[������ �2:��bзA��9P5�ݘb���@"��{�QTC/'ǚ�ĉ�\�M`�pE�����;���T����GNO��ӂ�WMɫ=�Wq��!�U6���}��˔�m5�V�Vx�����?�
W�ʕ���f�1%�b��sôw���j~�����;�N-��Z�ۻ�F�_�^���|U]]>�� �7�'+�1����غ���D~qII'�bT�^���{ܧ0d3C�	Z�%V���{/�o�ٳ>D�H�r�T���,elV"��>��$a����Z(\OOOKK' ��~�r)��Β�fBN��*��R��XQ��h��Ro��+�+��\:tamm!`���i�^�w�} Q�\�և�}΀��A�^��i�.��g���b�v�R�by��Y4�%�lE0�X����G�d�;����m��%?����W̑R�)�*��"�oox�������䪪���Y�U1�=�T3�X��ý��o;�A�s 갇2�2��I̍��A�
De�>,�"f��U�B�f��S���j��0�6��B�R[�1�-.t,|�?eDW:�b����U��έ�Z�z��N2��^�����{@)��}D�e͚%��W�%x� ���Xu��U)���GJ�` t�h+�K�"�zNa�W�y�@�����7Q�̯F/ '�h�,K�w�6��ro�֚m��j9�eŭW�9ݽ�ָ��Z�����T)�f�b:Pd��;���� ��P��ңV�:�'��>�y_
��H;������y���AC"��9�K��b�s}w�$�E�v���� �@�&&%�n�Ei��Z�vގ��*8�����M�������U�[��r=��<]�U��̥�얒���W�6�:���_��텂h3+���k`���rt�QLZ	�<֢�
�[{1'=��֘��?��R'&B%$�ɜ���n�O!��f���`;!�%׳zBlP!^� .�?���O���bh�s0��l�Qa<ɓ�)X{�ռ6�B�97��}�h�伛*�b���f��=j߼z%��-�Y���r}}]LD�[�=�����5gMYv����,} Q<<,o+���)�D5�MTcIi)2e8*89�����k�&�׊���Agi�ʲW���] f��W���u�-����|�;i�?�ȵ����O���%G|�76�){�VlEӒ��Eʼ:c�j'�5\�r�1�G.�&���V'7k#>�������x��[|E�d(P�o|�����A_�B�����+T����)�	Wˍ�˧��������!<� �R�i%Q���#׽!��f�w�T5O����8��l�H���}����K��:8��|]�������*y�DG��CS0arrr�ﺌ��)N��J�,U{PB|H�mf�����&E��Ez���rF�ѥ�oĵو�cf�Sb��1a:��`N���u�;��;������P�:����fBۧ���O�f%Yn�{�޿��xd�������*$�Ψ�BO�����=���T."��
�׸���LG�{�t���*3P���$�`pV]��s�]���0�˗u�B;��d�]�\(�{�6K�6s���-���5�f���kY�b�,� �ey�l��uvVK�G��:� �¿|y긹j6I�{nr��nטo�\^^^v�{W{����X��W�X�K^ޅ�
��- -�u�~N��|1�BBB����-ԧ.?��v.�+/:::�\ZZj�"D��俗|�4�#��t��X�N��)>钘��V�&�=p��:,���1E�A��7��ʉ�$4���ri	ٮ�ЮJ'�N��PHZz��NMc���P�q�v�)^9G�������R��F^B��OL�߇�"3������Q!X��j��v�눡|#!����g����4�����?C����5���/-jX��0N$=��M�{�PǀZ5�spa��|F�ِ�Ƿ���?*<�m���Y[[���~3v����*םP|�W�2נ�?c�{9=����n�X괧�)0I��������}�=ϑX;���������`Z�'�e����"�Jl�!�����<�K�X�=R�_�����Õ��|�:]\��/2��Kt&N���GG��bp��zTĸjn3l�5�����b&�¢=||
h��1$�W15W׌R�WqcR�Y#���3�>�v�L�0��`�闒�1�Mg்	��C��T�{�W*��ߟ|�d�`�Dr��Y�̸��>0�$���Ao���4M�<m �<�F�Yx`��'� %D,�R�������1�#����I�j�ֲ�+#s��f�K <�~͞#�勼N�A��04���~���j���D	ZvcZ��w�eo~>��C�K�bV&�r;Z Y�@5�ֽ ��P�盠z���z��is�Z��(ă��p�f��� g{;;5�=����&�e^ai�˸�UDH���-1H�No����*^�Q�Xx�X���ɮ�}AV�(�ޗy�\{?d�v���/�$8���z��'�ڒ�9**j&W88�Dl&��#>�2�{���VfO|̀�jhiu,ME/}�62ʇa���M�n���;ς�	@_+��@pq炓�� [Q��]R�1�U�^�NNzV��Ι��O�	3(]�N��X
h܃�n�����S�vf'���ho(����\�S}Œ����Χ�+���W\����2o���B�\�C�����܎F>�g�"G�յ��=7s0�5fB ��P�u�l(��M�XmKK�Z�F���} ��b���`�Zѳ���5�� ��_��z�%w�oq��qٕF�&;�!lQ7���ַC�V������	���K�����[�����~�ˇ����x���0R�W�3_���,����Ӆ��\�+1�#�"D�����`>���LjC$�YZ�	˧l7����$&�F{~p�MNN���r�Xzt���j6R�m��9�����T��ٓ%d��' s�n!Z���b\иw�֙39ӂ
�&�� ������e0��iii�K�Z�Kssm�Ly�]H��R��xH��y{�'��b`���na๠:����7�� �#Wc���K��B=��G!�8g�@�\F���T'=j^?�!��)��Jm�qG���5^�Qb���֣8��ք���ۜ޴�n>�`�+4"�L	+�K4�F�i<m��??��8@x�'�j���U	ߑ-�HF]���4�9x�_7I<p��Zi��\=�&==��N���};J�	��ydE��G[��i/{=`�,�o�\�{`m�E�Z�(�W����a�z����3	30�6yb�?h����]\L̬5�8�˛J� �}���� P|y`:���k�u��!>�Q�uϞ�X��G'g���$��0�C(��/��m��zw0�^���j�|L*�8�d'���2�p���?���0�U��.s\Z�=;�;�<1;77ݕF,�o6HMS�)���t˽r��C��4!�xBG.�����bE`u�(2E`)������~�G��hL��q"*�%a6VT��T��o��ך�le�$�D6±���9� 5�.���ևz;.q�Ĕ�M^��9�V ?������&/: �+��^�cvj�iMM� M��|��և�ӡ'_D����A�03�ܡ��@��H$i���3|�����@����C���~�Y:Mc�ޱ߳-����s���?�N���߷q�!QL�`��ʌB��1H	�G����!`[� �}]"���:	Eɹ���c����J`���逬Yߠ��������������q�+�G��ب�Hp��-��.W7�Be�7H�l(Ž����3��ʣ��Y�w���D�p����=#��SW{��~Te9X+�R��>+�X鬚Z$�[�++b42=+&����NWV��&�C��@�>~��~�fj�J�����7�(쟦)�?~ �F��qq ���u�=xp>g��ۯȾ���p��F��Fv���$����ɞΔ��Y)��x����щ��ݺ�R�l��g��_=+�X�:5��tV��^��а��m��(�Y- D*֚�*]�
�dW��*�*��Y=��������C�?&�D��*���-�
2
|�~��F� ]gZݷ���W��pU������;{V�6���:]/�z{��;ϲ)l���^K�fG髨��Z6f����#�����2��$i�#���1�f�܇0'�}�&�r	i�r�Ç�`���Z��D�_,�h��̙3E��Z��Yb�p�lL(�R�Уߪ7�`)��r_E
[%O��;�

[\^������ʜ��/~
؁	�P�p������[�I����]�é�1�DE���yN�� �O�
��<��H��?^v�M��uŎ(�;F졘[��fFF5��u�P?��������� ���N������?��S�G�Bq4����h�����ު�����1��JWQl�-�SQɑ�j���LKg$Οp��#$!�TH(��w�<��IX���#hi�Hr���藯ױ��cRѥ��M�������g �ݚ�_�ܽT�D����!Ӧ}���[� j�9����e8����>Xɼa��K��)d���jg�#{i�Ct���҂R��z��uz��sz���9WR�!���لh��Л�B�[�8
r;2��p���ل,qfxr,(���M ������!uZ`��h�;�i��KuEB_�D^��{�0KT���@��؞㙚����ю
qq�\�I�%&&�?�*<�W]�W?�?'"Է�*`?=]0` лp<�ւ�u%%�i
%ɖ+xl�|��''����v��7z�3%�lT	e#��*�N��l ��ӎ8~����*�;{�ZX$5<�����L��~��tu�QfJ$-	++^ ���@�J������\���`��T||���oN��8�PPKM�)� �2��	�l�WV��P���,�B8͉ͥC6����e��Vqj(�!l�/>ڂ��Zrm�+�r��ґ�����ʎ�
뽇+ݶ���!H����<G���S���0%Ƿ��ب>X�sB��t`6�e�B&tx���XOONJ-;�X��)IdJ��z�b�����*f�y��}m�O���7��ACV\��d�	�:߱5b��8 [�?_�,�ޒ�{�����2W�R�ck��V�l �D9y���I���\���L�d?M�&`Ĺ��4���JA9z��F��%�`i1�rtv6����TW��)c�ӽ����}$�%�@�k��y ș�U��� ˻���-c� 7*j�\�;V���Ԫ�
�Ð�����_6H���R��8#�"&h���9w,���>�yP`g��7��X[[��k���w;���[Y)���H�C�He�\@Nb�i�43��:��?�s�AC$����e��f�e8��È��`�Eμu����iG�і(�T��u.�����i�fck�&��fi�5��	�
�#�D�dڰ�����Z�	�����y;y�!���D�ʤP!���'����}|�������q�ҥK̓n��6]Z�I�����������=:�_H۽*%�#�����?}�]���^�5f
����uj��&F_(	�i�]r��e�צ�kK��h����#�6M��ț B��iժ2,��������-h�G��/��Z��:�A^�piX'��v��������>��Uy
kN��� Zpt�Se�F���	��u��%mٿ���m.S�2\A��������;@Ę�p��^^՜/|�*�����K�	ي��D�q}/�+{N(>��1E��-�_4(6�l:���v]�(��72*� ښ���iZ#�]��xW�dM�l��D<�fX�9ڳ�=U�/��N��3��\�ٮ���h�?�*�^�.��>rH(i��pQ�Bp���'�PS���2v|�	cK�*@V�>~DP�$�?"�&'_V�때��"ǆ�땳d8�8��>G���������8��WKHHp��= z@*z�	�b���ǎ"Lu��5��Q����,��Aw~�Zy��x]`�}�����};�㡊��$nlЉIK{�G�fU�x����|�E:��?���͛7�	I2���3H###ˢ<Ժ ���q�DɎ��˧���Q`@�~�x�1B�8������FO�s�p�^���w"�NFZ��e>VU��l4S@6�����1?�J��?��L���?�Tw�A�ς'C��
�|������{`�Y:k$R�Ģ���GV�!VwwD�������C/Oc�_���C�T	���:���{i�mN�fG�H�l]�1'ln�j��N0rM��u6�����f��1�{G^M�xIG���>!�BK(��w��o��g�N�<�����	$xp!'�F�^"o$$"r
_�Y=�������'��)�XOr�����`'�H#3~���U7&��\Q��z�'��>���ϋ�b����Y����#YԲ��i��⋠�u�u����^��������VUW=y�Ϡ8A�r����9YYV�����+�"�8���C�������yS�!���愝�לi�*f�vU�܊@�b8R��+�Y-���2A�ڟ�Xj�F����zpW�RX�����E6h��l��=�nڊT-`��|o�e��ez�/0�[�%%%�9��L���t���*���2�V������y-�IG�ť}�N�c�O�F������/��>_�|
-�_��А	�2!�22��=�	��n�=�mݍ�5(JQdU�.#����I�r�{�#�9�Σ�x~��	��,@d�ǤD��zZAN�3����������G�1ފ�2d���-���v����5r�u����MP�E~�Oډ�?
����N�#�݆������]p+%�X�,/�������TS�=M���
@p۰�q�EAU�g��&7�M^^>K����2�����_�,P��K:*T{1���Ç���)))q����5�������?=�p������	Tf?Ƚ3�_2
���hAr�QW����#�����ص����X��������Q����F`}`�<j���-������&{�XCSɚO�cT熉�y�[M�h f���Kƫ�w�� +�2����f�%�s���R�Z����(��SEqT�3A/D-��H�M1Z����r�u}�G|�"{��%u���gFbg���Gw����M�h������i�Z�n�ö��SL�?���|rz_Z�Ҳ��)hx7�Wy�`��Ƙ��##�N..�k-��Y�����/<褔+��7H�@H����=���LD���|vO�^�w�wy`f��q	��F���]Ȇ	9�w��-�rv�8�w2��,��QO��n�h��oҼd�6=Pb:D$��f��9$��$aA&L ���z��c��"����S}��.8�*-��j�-��LLV�Pl�������ޠ���<F��	�T��:uL�!Ï����g�f���V��j��,�m�7e;�i�F�333Kϙ�95�!wq9?�G��C* L� ^L�2���\���nD޹o�0r����*�@���;�{�3�:�b>�e�����ʀQ�ʨ	�޷s�w��0��d}Di� A��<E/�!�E�!p)!ezj
)Yd��>�m����q"�+����������g���9��uy�eぶ���?@VB��sz�6��L�t˚���G�]���A�L�u^�eĳT�{y�Y�^�mz���R6$�9��?N��6�|7���R6eYn�gw�NZ������M��@I�2G=�����>̌q�Z`13J����}X��S�>��mYl�6�.���ċ%�� s�����{o~��R`X���CYn��TQd��A�](6u����.{�h>*cg�=�J�{j�o��)G3W׌�o�VnRZ9���Ӽqe"�}7Mپ3�q���'���=�L�J5����;qh��o�k�|��	�������P�+�puՂ��^���6���*1�Ť�#{�����+�O�W��o��iqW�=�L%�A�y�b$��b!dupQ��v��{gԺ�.7�E��{ڝ��H6v,�Tȗ`�[����n�A��h��]�١q�j��w�pOZ?�$��g��^�[tC��a���}���69�n�������tx�DƔ����9�f�^�2|3��j��[��Q�<V��>��G(�2}��<����¢׆e�� �׍���~\��m������&w�f:w��]��{+�o߿_��{ �]��%}����S������|�V��2k�^��S���d���r�V��O�S�E�*������^iۯn����.��X}ek��=p����~j˧āCD�P��N��~ԡ�P�&��t�gO'����D[�ۯ=�hٽ�����45�O#xJ�tĊĖI�Ǐ��t��u��a��s`�5���7[�y���W������Q��Z�XWZ��Ӿx���0�!K��x�����|<=�����&��)��Yk�%r��%�q�Se�7E_}���HP=���Fߗ
��ӷEm��V�������I�b�#�y�4�Cw���o/�X�4�R*i�ׁ�;��Y��H��ȧ$Yn�9R�5Y���^J���o��3g��5�DFvh��M����15�Z�?��|�c�m�� ���soǷQMee�>[}�MBr�f�&>^o��{[G�w����t��$����ނ'11qt�ǹ�v>�۷;���)��yxZ��T�[���{v�7��J��貀�鎃fBǋ��zS�<j3�l�}W��%z4�va��/��:�7��O^y��5LȚa��^�?��|���TOXx����p��p�7�inN���$w���|ģ���4��54��1)�~���ӡ����C�^�tH1o�r~G��i��<f�r���7Y�H��gEv�E�n_lcL�ZJ�����$�n{�|n;���ܼi��%vq�#{��~78OH���q{o�/�H<�5��td�����W��_3��~���}�Q��	3&�eY�5�~�$�8�|��	��k~���J〟9��m���UEDc����W���������?�T�-a&4s)V6�#�7t�5LgЬP���&-��f���֊=)�бG-�?�<��3���Y1(��n����m������e�
�p�r��s�'��=<8�3(&33��������K�z�||�C�,�q��س�|."�R3�O��9~���QX�Ya�'<M��Oc����g�,g�;��Jw�9gn);38x�V�M�p�����~����j�)��,C3�n��1�$�3#_'6Ϭ��&��֮y)O�N���@V�՟F��b� =�~� ;�^�cn�H�:C�6(`��������� �/�B��n��((:���RC�C�Bm�Z����b&�юU&%��sñ*Ԥd�Jen�#�ee�-,�k����>�����x��sٯ��{�2������y�u^>�d�f�
�:	-���"��E�
�b���E.nn���ZCG�������u,�����lN���BB�,�?"�I���Q$�:�WI��^�ɖ��s䟉|~���w���.�
��v�w�i�w»�ˑ�1��#�N�(g��uƈ�m��	HH�x�RK�ƨܼY��}
,#���o/������g�og���A��6��v�rMH���W�Ep>�*RY~\��>��CrRz�"�a������No�J0H�hCv�Ԩ)�yY٦�an���g�޽�����fY昹�Z*˰�Z��(&���y?�y�@�:��Z |��Q�&1��|RGA�~�p����Z����'��@.����P���N���@/��b���r+=s���@��������x��]�R��x0�{,e��V���9A�Ӏ���Gz�{-1�����*��V�JZ��������?�1�6(����x��ϥy�F���/� ���;��0�fBUR'�VEaG��,�}���I��w����E4���D�_�hI�La�ȜY�"��m���u36���ϐvXŧ��4��{�b��#7�;���?�7ND�k��hjI&W���-�ѽ��[���I��	�l��K���f2x��]�y�4��K����Z_bL]��=��1��dxee�8۵0lic/�\�1�!_�^�o&ًmmO�4�l.�!�q��:,#[�����ޞ��R��(���܏�.6�c ���n�U�LJ~����œ/�ki�ڞ���Fj��Z܊k�ԗ�xrS)�jRx�36�Ѹ鷵���nxj��U�54�v�%�/��Tn�Fe��ӗ�(��\���7��ך]/Կ�`1��u�X����w�o�~|��&�����k ��ॎO��О�yp]�qK	hT�O�ߓ�\��s�2���^X𙙥\�yb�B���ƈs���G�F��E���et[c�/K�=w���1Gr}�H��>�V�����S=�p��"����	��cimt٢̽,�U���B��k�L�������a{��������"x� �*�t^$m�y�9~2*��SCj� 	ʅ�~�
G1@"��uޭ���?''�!��mL������i�������q�4�������5x���z"d�A����q��C��Y��ߍ[�T	޾����޸Al�  ��!��n�̰T�j���HLy0p���˞���u ��eއ������r��8�x�C-d��H]t�a��fc�! �/V}3g��SH�y�c>9��2��ޛ5n��}w��7�
�jHV�w\|A=���s���>W��n@����3lwo�4"�n����}��Q<��ɓ���o[;;��k&���F�[�bk������W���~=�eK��6��Na���&pvu�����F���^Ʊ�����+Jm�}m���!T�qlᮣ#G��MF����Ǻ�}?m��t^�_�A��!���Ioh�8p8Vz�ܛ^_�x�78�����h7��$�'��?A���P��>�<���-��we�%�bv�"��
�������~�i�6�z�잣�A/Gᤎ;ƾ��t��%_m��+��,��|7,w���F�ł��r�ذf������ě���1%8�SJ���]��--��#��0�)+;��y fP��tP%��oa�g����ҊG��4X�n�ڻ�����.��T��Afp���U&���W�PT�7�t*���fW�f�W��ܛgW���@8������	�,m�E�苇;ǟ?� �me̪��𫍛���I"�ˡC�����6MO\\Kmn{��������ya&%��:"{�����|��B�>	_��;0�t��Y^���L)�T&~ϣ:z���D�\��3.7,�g;~�}���mR���Ǘ��h�f74�)����o���N��P~��nΡMsҿ��b��{�,J�&c�ڄ9H�#�8��0�2#Y�?�?����y?|H��ᘻ�m-�Z�@;�IӔy����;n�ftE���4��ue���q�{�oѤ�r�\ �K��Y��@�f�P�26O޿�x��|'�	OП�]]�2\O���z\���{�贸v���H�!��u�H:��y���+@u�	_��>P�9e�O��s����/���	V�3Au���+��|D����j�<��,�O���fЭ��)���ƬE�06ߕ�t�2ɷ>Jr����v$y[J,M���.r��k��A�ϟ����ʮJ�D�k��T�P�+�Q�c����>H�U��~�@o{�FG��eT�����3/y��t�3��u>}�.�s!�����.g��۷�G��0+>ZvG�����4�����xr�Pv�p�~P �Y�o!V��q��9~e�¢C�l.5d�=���U�l��⚬j.��'�;�т٦��5 ć�K�|�y���_(1�8z��;g3�s���(�G{y����(3,V���l�&��\q�~)��6�-*�� �<ls6*M���xƳ9���z*��:��K�ΰ3Y,���_�fH��py�}����>�<��	W]�������:��F�֎0���#�i��}�^erc�f�V���m�Ko'ڮ���؂#�y�H2p��z���^9�y4�x�ax���W�%u��R�}4;{闇1]\����33�ۍ�Y�[�ۭӷn*�?�~yY�*�2zW��"Χ:�A����$Z�n�h�wc�_���y���$nA�0��ks�;�NI �C�ɦ��޽{��A� ������S I�ըy�ϻ"���d�����v����y0�$���_M|]�E	,t�n�?�afBa�t�dOT���c�c�9�t"Z:jvVW���:�2%���a��1��n���X4��9�-��i�j���;l��QTt�e��\�X�h����q1���;O�w��"4��z���!w���4��Ю3gΰ�4���b%@����h{�@�&�8�}��,9t��aө{�7����z.�eq
?�y�e���x�����h$"�5D�	���D�����cbN(�����V��!�	c/x�Tx/$�������S�XE3!BʲߦZ�":��C<�c�<�u���>���2�yi�*ZV{��F����ҡj�����)��s Mi'/Yݿ��Q�O�!�W��jI��4[!�׭�?�������W	edeoB:���HBfFd�ʖ�Yd��|#�!��:I�W���������o���ܼ���z>�������z���a�%�B >�۲����P�s� �,� !<���6�].H�/�a-���D?&���t�$'#�@��X;8���+�������������թgOk���LM��ξV��ә�t*�����ވ�~w4XY����f0�S&o�C=;WV�|�����n݂b����fnn��^�3;3��Һdh3h��8hd�U��z ��0@Ɖ��`���++Hk�]�mo�m�(��B��R�o�v�ѣ9���=�B���qh������S�z�iJ.g���}� U�J?ԣo����tV343���~L%�thH_�����f���Q����C�#uѱu�;�`0~EV���{'��~[�2ַߤi
�/�֌Y:sPZA�Ze�4���x
 8}�+�G��_Q�uw�8nke�=����/w5+���X�u�ӕ5��9V����rJ�
d��_'�re�KH���$����f� 7�bx[0�o��X�m��=_��܇Ů��o�w�z{*��X�D@u����#诤:�ܔ	z��a�NK9@R��}V�"��M"��K��'�P�_q��J��&�x)$-��U��+3W���'q�j���9��a�3�]� '����g�ɕޙq��r�{�j`c�M��Ж�`�G�NWrWj�#�i��\*!!��@s6���==�GF�o�U�&]]��L_���G�3��@%�0��Ě��b�,p���i��{�Er�l��E�R��II?�[zWS��e@�4�(6��I�8R��$�?�Er��ru(W	2������Z�}Qq�`���Q���!��7(�P�*�ŴM���ݮև�z�G�1��Ύ?	�.G��!�1�_�O,��଴>Fs�H�� �C%���ɱ��)���2��,��� ?>X���a����;��������i�N�8@��v-+s����]�����5��ۍ�Vo������~Ŝ�Jӗ/ܴ�r�q]*��˼���""�k���P����n�EtN�⡖�`��}����R���?� Ӡs�)R^�>9��C?�Һ'D"1������m�MNe^�&�A�!�����ӓH:�x����Պ�ʮG�4jQ�3M�^��+�6L\�Z��w��A�k������� ��c��}�r>>[?�ǂx�n�ä{ֺģآ���@(�l3(���1�� M�M�|������Z9+�T���1?���[l�j�Uhϡ�L�Y�h.�<��{�I��'NU(�Nr���X;���%%E0YР'����J�/Ts����Q��5���8G�I����B!���({�ʡ���%��ALq�5rC�a��T�5�&�0��A����G��"�o���ᰥ(�k�1o��GoK<�L�Fw�8�n���\�%"ϵ��ԩ����mw߁e��l�!�0�z��ήT��gB&:3D>>����oz	&�g��BCgr�\'	n�TgQUE�֧��2F5���CN�葶7��&�̖WP@���P�d%+��Dx
���z�����R�;��{��ȯ��Fړ��АL��̮G{��z/

�n����om�����C�� ��͍��d)�Q ����r���lePP T��fQ�<�v���)����n�L��p���c��&�W:	a��n�6(w���"���U�ԭ��ͼNL��Z�=����k��
�+5=;��&姅��_z�D��Fcc���,����3���47W��]��NQ���i�&���KL>��i�9��o�iOOv8ԞԠ�/x��Ƃ�`�1�c��j�i�ő�w�~`�@��Q�N[��}��z�8�v֓=Q�����
�EA�'�pm�$edex���f��H,A�Z�ܸ���s ʟ�ΐ�N��#�:�n���}�'�����JJ��[����5m}���i~���~SSww�۷��~C~�SɕX'=`�Q��ï��U{�������>�뇠�d�����re�ژ�$�&4T�2���oj:ALӥ�<����c��!i�Ew�z�%��g3��Amm׵�[�Œ�x�d�5r^ۀ_J�K	9����=���R{'�������5n�<G����+s�Lu_9��wx*�
wG^^^XT�d�;���C߀:��E��u����.��#-��3�c5x�=��}9!a����
��ָL`j�M��<%�ׯ_��tjA0�uo_nϪ��Zh���f�#�񀋋�u=�x�wM*��%z3�ޏ ,S���߬Ӭ��*�KIO/(��C�,�p�P�y⌜Q�VO��M+�vVQ��_W�}�4z=""⿁hC�@)111�B��k�!G��9���.*ڀ�	���*� U��Qg<��F�j��o���n���X�w������Q����!A�0�߿�(�[�z�=O\�p�m�!M3J�S�� P�%_F��[/gJ����r��w��hv�}xH޽�L�!����78����cܜ����K���!%
x��u@߼��Ȫ�bpp�I��c7�i[��";��J�J��p�~�qe�s���t0�]����hy�,E*��_2���'Cg�������#u�����;��Z��3�N�H���٥�9��6�$�I�2Pdsϑ�RB�QE�R�7�����b��Ĵ[���L�l׀�ba�x���u���Z����,F�\�|5w�E��ő �_0k '�%��I@nu��� H����SS�2�%��[�Y8�|J������n��q��j$~�n�/�w���j?u�1��NZ���(o�U
���ׯۜ�;j��N%''�ӑR��#<�0��f��#;f�뛍h�M��ؔnUt�lgn��,��f�?޶��j_<%�D~�>8O�[����iJ�~/Ýә�������[�3��g��3@�v���'�|�B6��hÖ)'�����������b�٠HǝN��yҟ�����,��w��x��2;ղ�{Ɩ�Tz�����/��i_����ĉ<t�UKo,�`��h0���?Y�N�0i���6p�@�M޸��BT�����뢂�<ؽ�V@,�IE���V�j9B2rrS''����+��**�>�Ds`/��'B��&b�Iy��H�
����Éd|8��$O�(�����w�.P�CQ	ķo�Z�L�K?ϯ�<�'��^��Q317gM���Qm��6��JΚC�����~h�(��H�W2�x�@�� ݫ��� '��ۤ�	�A(�$'�t��֟����9�R�x^���6H�?�00��0�!�(��?�{{�.���UU'?On�Y�Y��蘵
�ڊ1���.:��gUqG�-OQ0q��g~��C{���kQƣ�R��(v�e��*�K�Ǐ�.ɼ����)���#��e)
9v�u�I��EJL���6+�>#g��#""J��PZp�<w�*\��ל�����erP�r1ErQ�J:Y��X!饜�*��>9�UQ��M�=<�Z�̫���� ^4�D�u�e)���gdp�'�L�L�"E��f�~Sܺ|�������*�?�
'��xv�d��|ae���0�\+�Q��<�/��E{\/c,�F�WԔ�7$�E��a�I���@|k��qs0��D=������{�	"��w��l.�KSQ��Cm���K��b�v)�5\��{b��z��靝WIw���=z�?8�X~�Z�8��@��"�'/'W� g�٨H?Aֿj�o�OT6a�Pd��-�/��䱛"Lv�ަ�������]C�FC2���P�f��*R���K<r�q�7������.�m�[W ���P�O�^��>>�,Y�f�����g�I����~f��I#D�A���8\^�t��Om��`�D�Ɔ�-w~�Bssw!aa��"�o��8��%R�BB���N���G��F5�k���Y�5�=��JJ�<~e!��
p��j�a��	�Y���_�6⏸T�^DTk�0������4��/#)��cU��E����122���ʽ������Ķ���Pu�d>$�������0c�3-�P4�3A�J��䖷�׎�����^��T"۔Z�l�RR���V��yc��o���_K�K3PQ*Q�I��g�4v��u��^ryj��uF�٫=�L���F%��ؚĳ�'�#�ﮪy\\&�����Vc������o��_�������s_BZ�etTP�bָ��� Ț�M	��q��!3�)i��\y�O���d�L�\��z�ӂ@i��ݫiBr���2�&�Zװ��jkq�81 _�B��5C�㿝�#,��x�7�H�`�T���?O�ò�(�>���ϺT�4B�HE�i+Mt}�a��tI��IIo�ּ
��-=�~9��_O����`�f���z�n�߇�BC�6%���s&wL���k�NhV	s�Bx��Urr0���ZZ���6ށ1jn���&�r�8�/��{��{_?sTo�����<���#��
׳&"�Y�YyA�s���R�K���~o���h���|-	z�]T���9�>jjj�jjN4	!R�˓U_�*HBx�b�[����'��2�i��pӅ�dM8��a��;����ij	�'7�F+=�43���&����dEN�=�_���b��T R�H�g��xm�}s��=#W���P6�Mn��p�ۖɕ����Zڈ�/
C�8��y��𡰄�EA�Q�DWV��ŬF&?���͝�RX �<<|C�5��g��3(K]c2߻�+��ݎ��l��v��ݔbk�����Sl��{��鿺J(.|�o~���ޞ�-:7�1�b@K��󒷽��t<�N�j��?/,�H����i�g���q����pV0h��j��H{s��Y���uI��⫢/�ZO�C�_�D��mF<�op֞��PH�� �u�GR,@���Y_-/��,U������8!�}**�i�7���w��d�Z�����������3��753�y?�M\��c���n��}�Qׯ#�l�� ���e�G�O��/ܚ��m�iz�\K �[*x}l}q��D��5"Г�����xx`u��F�c���f�Agu9J0�f��h(��ޤD�0E����P�eQ�w�����l��oo�����0���R�mW��kN՟��%
i;)�%�쯎�#ћj��^U��#橋o ��qI������.���iC�az�����U����[���tD	9FfQ܍��j}0
{�հ�O/;�84v��adѭy�Ԑ~�,V���f��ǠN��&6}�b�@��ɤ�-|�Z��`O5x[𧪻�E`L~��FDF�����5�.O��E	b	��� A�� )�����ڜ��~��J0�ˋ�����*28<�z�3z}]��Z48V�2֒�ΝM*2"�^��i]cc�kT�G;��K���_{�Z��N��Z树^Xڷ�G>�E��R]�)k��?�U>T%�_u|$S@sae�6_���f�ձ���;��G�ѥ���BBB$zuk�CdM7 �p8M���pӀ!8Az�"at+�t�A#;;�X@'M�����5&?��Űuc��Y�<a����maL�PJ�Sa����s�r�k��'�ĎTz�'�?�<N�+VZD$��n���r����1/��dj�<sڐ��l��a��iM%w
*���a�݆�&���[�!I�8X(L-,���$����o>2�04\�ܶ���-cX��)��?��H"��o�{my�~��izU�|���k׆Xx��	e?����؋o2�.}�	TxӉ��A��0�$)�@���h�e횅�����D�"liD��hO�����3~�彈bS��߹s�$xA�2=5�MJQ�>��Ī�&C�B���W�
k�Y���ۭ�n�չ�b�}@���~1d��?����BO�}b"&���yo�,mTT��iWrZaa�И����g�f�^�l�E
;+��@:N���5��H�S�P�oݯ��#����c�t���+���,���<D���U�^nؔ|�w[1�yv����빹|@�Ǔ��� ]�p*n�:�UG-,����_{��Ɨ�.\�1G��'��g0ۓv~�74;�/��]�{�$�)�LE߫���ZC���"�#9H��7��W˻i {�d�7�5�v�w�d}�@��L�T�O��$%%��'��<h�?��-�~$��X3&�'��-����& :_k�訓�Y׸y��_�J�͕Z#w~Ʈ^BY��vui@i�X��c�t����Z�)R~R�}~p��X��P>==�@%����6L�̃��⡶�fU��S��0���h'wN/o	'C=T�}�ܔaÍi�Y�#���w�Vn[<���/���˽����V������!��6qq̏�������1�OU���Pf� <���]OIy�)�>V��k���11T(��ё\���G������m�g�n&�R'Xfh	�\[�E�Ʋa~�&m���f,a gDDD���:�@�B�1>9V�{R�������\��i��6����Z�),��9r0�&$��	͚ ��KQ��}���������,$��"�z�֙���NwD	N�qE0.*�b%��0ٚ=!�4�ޟ��qt���!���Ujj 
[�b2����7���}�#�ݜ��f�++�
�z���א-~J9��GdYY�IRmӫRR7$S���C��>����N�`����j�iT�NIi��yU8hVr;��f_�H�!���[g�R�S�QeJ�w�CP�r���v֋�n�K�
W�>�m�c]�4��iҞ�\�'�^��_����7 �f�|�=_��c2&^��-���TUUA�L��Ry����op<�j���ڜ�2E��� ru������m;;����0��#�h�	J�*�)j�i��J}�G����7�-e+��;�}��suk;�]}���� &�a��Y�-�� ������C��]5$6L�l3+�� �Δ��T/!`6�7�)pq~># D��f�]���
ٱ�##`�`T~�@[,�VLݳ"`��� ݛVy�0�ys(A(,"��%��E�Z�h��T�B�Fy�X48J�Vő�\����M1l�{1��wE�2ńU�4^��XI�9
?՟��J͹i��r��/]��&u�{����J���A��ƺ�[�0�:�i��� ���L��o⽺ T�**����L.g&����8�7�35o���
���ne��0�'G��/H��)EZ�����1�(̤��*��Bd'���%d�$@���Y���1� �[�}�E:&��hB�L~e\�8��pexE�LBa���!�0P�Q���Fk�fO��~�C��sΝ��5��?[x�}a�""�)a��@x_�����p>��)Wד�D2&��'aP�`e���r��Rr�����Prۃ+BdYr���3����ԡW��U$x�7o3�=|L k:�*��EV�0��h�У��}3��,l�į���N�?����[��"��'�:{N.�$K�0v5��@���8͇��N����^kvC����Ca^��Ҍ���%�%�7�||�ݥ=[\�����+n�������8A"p����)(Î)'S2pM/��K�7eh	�ZH���:£�2>΁`��ǝ��Ut�HG6���r����ֲ��A�"˃tt�Bt�R������V�H>×ܞ2��rRc�[^��־��7��S<�fL���a��g�O�/��v7\^ZV���R�7��J�7L,��hl1�&���,ٯ���DȡB�%7�Bj�}�Kd]���u⑾84ױ����O`�a�˻'*�f��
�y���lk������3/��Iyo1�H�QR]���$t�8�Gcd���I ���r����9�7$3��w����Xv��S�`����;*�3���w(��p��"���o"��2d@��5z!����8o��n�D��@����i�26��w�g����yWU��V�'���%��`�N�Ğ�3ɓ����E�,��ڟ��|��L){��{�%� H��f�s�-c�n��=��t�����5���k�VY�`��C9^KM�3sq�%�U�־L6٤��V�Z\��̴�u���޹g�z�n=/�?���1�긿9*�օ��:.��1	a���p)
���TW�E�b,�9xӒ��༏�ET�G1��>7X���-���0�����ݖ�8s|���Q�)�`�(���-�|�mz�EYXY�p?����A50P����\���N�#ǲ����說�������]�!'kzt�2W��9����;���ڜȈ����BQ��['N������Ρ(����&�'���$k@� :��rP��Ʀ@!���s�I�JP�i~}�H3_D�ךۯ6�P���SE��J&X�[L��z~U,�)`	Tb����&�L�̀	m3�,ņв]jņA�Q����f���<fܯ4��V�Ūh��*'L��TL�k>7[���ih�w2E���j�$��6Y�	�7v,���p�{�����_uuQZaM�k�!��SNFq
<�w�=G,z��B���7ksČ������rmꇐ����Z��?	b��% �Pd=es�G�K����������H�U6�R��,\s5�
�Mlө��/S��/��lū,��a(���TK�*�Qة�*S��]��)xWR���6O���>8���J_���fY�Nv��f�cӬ*��M�s�K��iO���щ��x��0G+K	��@�j[ �.�U����ﶴ.�����ih#q��O��"���ϻ����s{�G�w��B��1�9����O9��%������>��Bl��8�M�[�������f�?�wo�Bp��_n�>�fh�.�kH��KD+(���W�sNUM�|7h� �8Y���*�U���R��WB<�m$Y���q�������?9��ҲxC���8�@���j�ӑ��A"?�1%���9NEjo�x�2��a$�7";��mٲ.$b�XH+ҹ��3aq���H�sT�iݓ�D���h����l	p�m�,����^QY������8�T�+�2T���������� �[�8#�<�g}B��#�h�����
�����}]�����Z����+Sɩ{� F&'i�v�]R��?�U���������Г�� ΰ�:Q�|��gqq�,ll�B]���О�ɬ�����Y��{6m�KNNn���7;H���ӈsa�"�X�X�8[W��\%�QV�$�x�c�r� ͅ<��U�k��'�D�6�o����!��s������A�<�Pup�(.ʹ��L���P��͏SDP�Z��К�}�I�#�O�s��_�z�O�|��e�e�VI$�{}�.�<�2�I�p<����{ך[
K	��W��`���L�������(eS���qZW?Q�GZ��%0d�F_W|��/ ���J���/��fWa.��뾱r�kt���ĺ'�R�S�|�VW�P�c�e?��7+��IY���,�LJ.����PE��!�~`P˽�������P���n^E>��bᑑ�R>����ݍϑ�'k�!��4;+�U3�/�	,;1aJp�y$?p٩��+��gv.:���� |1;�i�y(O�I���#������|-�XH/6�H����(�y���|^y��J���ᚡ�����N��Յ/.��A$�#��W�)	�vtI�yC� W�f�jО\]'	n��{�=���[����p��ӭ#5�Tћ��ڨ78F)��f���w�&�(2��4�^sO�ܟq�w�`��i���5�Gv�H��4��TWW��(˧�໕�*�iB����>Mf	��F��o�dJ��9����;Z��/��d��Xk�6#��/,�K��!���w�1E��fQ�dA#&�#Z)�����ץ�Ɇ�NJ�~�8�4����\L�{�����4 <2�;��F	�p����җ���qy�G�|\U5J��ob��h��%
��d``xn�ğx��M��9@!�Ӟ�W񺁠8q����@MY���kj��~��{|���aw�͊�Kv�s���2�/��P~5y�:����2�'�8n<�#|E��#�����󏍇��T�a]+#օ��\��[�z��K�ꍳ�ڤ[��f�ÌoX��;���$�U�?�9��V��yu�G��}��u(r�R���{>�2�ݿS#���=��4)g�3�̦�a�=%�������[R�o_��okm�t�D@������ͦ�4�k��榦��2u1�*4���%����_��2�4�����~{$��B�;?(D#��i]��\L��������㓧c
~Q�x�U����"��nP���9;*�~�Q��N��!�����V��ˤ,�։���Ndiha�/��~�Q.��G�X_{��Rbv��"�뗘�7e�>s4&'�� 5	��%>74�"c��n��y��K<n�]^�k����\�еk��X��V��%p�H�Pu���s�L��ڻ\�W��6S��+F��MSH#����e�j.%Y���%R��dr/��_����
��Q[W]�˳��YH�6!���$,	���-Rl&?�g�wԁ:�WGQ32Z�{����w�[����ǀ_�Uv�33��d�ls�j�
_��_)�b��.)�K��]؞ק��9Ԩ�1y����f3]}}d�LD��S�֛���;9�+e��\}�"��tpp���'Z�t<��`w�#�tz����|�bz�h�v��A��%8���c0�]	)�r6�u�`hy���T�A��pJ�� �|ᙯ�Ț\����aIXq����	�↛;~�ylс�^�ecg7uw�mͣ��
<yG���5�h3Ҡ�S.��&&&�01���a�N]�����J�{��=�B�0.���U���-?����meo��%6�7'+Y�Vn��Z�Ą~B�y�Ӻ���ǯcbR*�~zzv�D�T������|����  ({~'8�W"U�{��q �BX/ �)ϭwȮD���(���7jjj%ee#;�=n@�X�渋Qu�r�HI�!��W��ʨq��X��gώ)t�
Z��F�W&��^�t����V���� �S�Xs���%�*p�n�%Oת�Ɖ�(�j&R��0o00/:h�k���;�o+�!�V]�ٌ��,��=$Ğ'���E޴��P����+�����3U�;�L����)���4��PUV�ΙB����&��G6ҽ�
���F�bH�F����W�������D��_������Y&�=�-�@D�YkU�F����c-ܡ���x0��r��b;��#��}Vw<�(�`� ٶR�J�X��������Urr�k^~��i�)v�H�<k�Dl��O{jM���U#�~�:U�������m�����d����w���,�?�"�(��+6碨
:�!���~s��b�����I�����Y\k�����Β��RR�����Ƴq�+����^2f+-��{�URۃ+W��9eՀ���#�h�V"�B�ND���IY��;=�	GB�����aqQ�f����E�~ݳ��J���R]Bc�d��\(��~`�Zf�L[��N����^`���ž�a�\�+[�ω&c����@ϟ?/��跢���p�U�V�d���2W��m�Bs=��.���2�(�z50?�<�桴1o\KK���G	t��S�1�+f���z��-�����C�%##^�d�ݒ����� d�ܮ��L�H������X!��)��:��i��{UZ940z��KetO��pŀm�\u]��6n�Qo��Y�����'V�;P��[+.h��\�eVƖ�5��$X��:9��9��o��wٲ0�T�Q���*b������ܯ����N����IG@.�����<0�̭Bdo@x�sʾ�fB�][����L�X��t���>�6I�Ut+�����5U�!���~��[�`�_|��AKE�r�� Pm�U�᭣
�G����o��ZÔ����OB+�J����M"Yt�l��%w�T�A$������LD�f���A�)��gl��)�*<������RʕLL^�?5�	��t�MRjj$���(�P������N�:��201�7M���4]�e�K�Zj�� �R��tc�->��<S��LyK���I����,H]���"�U���v��N��T�Q���4u8��N(���5���y㽟�Bn���d�x�����M���y�����6�>�~��`E�������ӌp�	�������>�:M���_���i\Z�b`O�9]ӽ��3�~�A�9R��W<}>x��Lक़�4�݀`��>2G��h�JY��i<><�`Y/>{��ԓ�I:6�=�0�����G:Y{&��9�|ؿ��A�wK�L�����{7��zV�uN����K�ld��7�9kw����#p��!�4���ء�%OO��GN�/Zq�j����a�1�B������z�� =������{_C�����4�>�2�����AI�Y\|�ך����+��W�[���O�[0^V�98R��52e��m�ኩ���`0�!�u��,�����Y%Ţ��dM[�G�k�G������F���s�t�{�&!�J�g~�FBJ
o�/kЖ|�`aUj�ˍ��������p�����^��?�֢�˹;������@a��w�o���0��K�d�t��G��D%J#_*¼Xҁ��e�Z��*wzg���sK�Z�+:KC����:}���c��C��8�h��|-j`;Wz�R���])$$'�2���LS\�ڭ��ëN�J�WY��3IC���+�{o��Vfse&ɉ2ٸ�G� s?檃��s�i%���)�>��:����/�{k�$99YHE�Q�0<����|09{�R6���9��s|#�-�t���DT�����Y�X2��mB8E� ^PL��?#x�rq�2X����c��*�O�Zy�۫1�$�����ln�9=?���2KG���%��I�G-E1�����m�� �X����t��Nw��T�kkٿ4	�����
���`̬f��|�=q"H��%
$@�-4Kُ�9g;�wt f��S���2m��[:@���7E�a�3�;����&W~�.Z��ҋ�x������ Y���_� ��>5#I_���o ��x�9
�_&�/���mtO�2�L �	*w��U5jT�%؋�J�b)��(s�8}=���}M͵���Y$:KWVN����^Q�A^��g� �0�(��7�`"/'ssW>O���e������B��Z^�>�|���,3ٛ�Ib�++`q�.E�	����v�<���9Y���E��9'@G
7Mؘ@�	�	���}�;/�@5�����>��չ��L�֔�\0<�"NB^�PMqT.�����o�[B���U22;��Vp龍v�B=�.�;N��,,T�l6]H���\�,���%w�������9}�4�;$��K_�&q�x�D9VRQfuM���[0�Ohl��+�11���
G9޸����JJ���/䢻�9]��$�y�(CK���~�.�P�?-F~u
�;5U-1ND[N�1�Ի���15�_B*�$E��A�W9Of}+�[�LML��x�IoGEG#ۊIy���ee�	֛n�]�J�#l>x�#l�2����e�����j�N5#�b�}�P 1`����D�
�<Ea)	���d)�
�$/9¸x=��n�?v��[q6��jlu����
Nzu��-������&I-~W2��[��((Ƹ3u���J30א�U��>wf�KR�9����9�0�(��ԕ+�$�M	s*�O?~�fv=�jU�(����E�$]c�[(:�'�\�F�οS��T�2���<}u
-�R��[C�=u������㩚�A��wO�޿�������R0�]�kdg�?&|kD��K |�3�z����ۨ��~��m� ��(���
˼���F�ˉ�g�����i�}�����S�
ى�"Y�ˣ��ߓ?�Df�����z;�rUG�.0�����jt�?X:�Lڭq��˝����b�*��C�Ρ��NG܄�iP���=�����>��k�֐�ly ?�|����L�+�~;T�lj5f�o��Ö|�X_b����q�����iU�}W��d`����upW��p�몴�Zj��-�~�ڊ�7��-Av�~�zE�b/$K�F�V�����ΐ��^*�'�Tdv+���p��ޘ��N@�=o..d�0 �+{d���}������DG΍���ͭ�uT
&V&o�Ӆ���^�P�&�����P{���Z݋�9����uv^ս_�W�p}a�`��������b̋c���^��ddff&�h�0�0��ں���m�J�\O
b^�\JBf�"*)),��&�I9��T�����v#4M+�� ����,��M���1�ŗUh���+Mi7y��vL�́:U�K
P�+����a����j��D�tiְq�J!d�{҉�Z����uk��BH�ޛ�p����hv�V�����.����!�^s1��#j�wpITelJ����|�L@&?8�2����C~ Vk�Ό;U����;��HzR�=�Pҭ�}�w�:j}]�'��l�0j(H�11C	�j�	Pqkj�J����{�3�'?ٻ�����˴�y���徛�k��%��{�%���_���P��m��M������n�3N�N!���C�.=�����q_�T���O˃i6�p��s?~;]�{�R�������',N�~?ZC�9ȴ��Lx������{9i�Du��K\��.HM~�a0�OF葵�[2���0�f�k_�� ��F�MKq[HX�X�B�fI���ْ�� �0R���Ȏ#��#��O;�ږ'�������_ݝ�ZF��ji7��L�,�?�������t��*��>opӳ�fKl�I�)��f�����^EX��	d��NPu��f�
�5?'@�~���'8
s�,E�ݠ�[k�E���z���S/����z��s��pRB����i׽����߃6Y��!���C/;Z_��%�X6�OQ��OQE�wģ8�"U�I�t���f�:|��g������g$�n�AY(}���@�P��m�ߢg&���Z�-:y2���aۃ�yYC��3lR�޿���V_?��^�r�c6�2�G����H{G_Z���D,q�UXb���'��[�^����hkʨr��(kk[�B�+$�Z��Ϟ2���ݒw�Hc/���]�M��l��p��$�=kGj�Uy:.��i������V5`?��ӀT3+	1+yz7>Cnf���J�uE����؃��֡�v�J����;�<_�}�-���kk���-�\��<	;��Ɓ]Oפ��x���}G��.OI82�D�{�I�#8Ů�k�Y �U�����R5�g���-�w,��0!'
==.#����	_�妺֨�GTU=	��m�8�l�?l0�b�C����g���.�����|*����J0�l�`")�}%i��ݽh�+&e��"!2��&!2��c�}�ID"*�&uz[�;c�K%��ȋ�VSI��5�P>���Eޞz�ڸ���ޱS/x���[�+���x�ض7|���X�I2uEfaĆk������raaa��9��7{�P����<0�{�sB�6�ԕZ�ʣ��
;s���i4����݀O��%`�~�Ђ�D�L�[�X����:��1�e�K��Ho�
��@!�zټ͊�σ�L�)�O|��:�o��;z{?1$��� ���QH�gĳnF��Ֆ����z�1��)������\��v�C3�Q�ìˉT
���T���z���Q�Z]��^����K��^�QB�q����v\1v��|�q0����%+#W���2�ӑ�M�'�!o<��XH�c�; @�?�"�,jbcC�l�q�=/��%o�v��R�Z[S.��:i�I<�\8�st�>�f�+6��'uk�~�"�7�d����WiR`�9
Uq�n'FK`k�uL*�-��[4=�9z�����iik ��p��w��DT�,.|Xoȳ�VVQ1�j0�LmY\;}R���Jp���	��̈t����\�]�B� �o���۔��Xe��/3�Zn�\�������~{
���gq�6]�u9�$�3������7���8� �7*���Iz������Wii%C���xh��녪PRR�:�b���<��",$Ͻ��c��࿷�֒��]�)v�M���L�M�>kv�����[k��K`�<���l.�<��q@�$������%c����yQUn�&�9���?
c����hK��?z9�@#���:���Y��[��2쳰M"��89�4���5���	@��ĘӞ�.�&K���n��.�R����݀V��F�޵B���Z+��WR�T{�n5'���H�n����ӂ�'
*]&��o:�1�4D��ol�ܓ_����\X�
؂<*yK�+sy0D�P���hf|؎΋]υ�O"������E��4
�G�M�`�"o��4~�<m�𻶥��&c<rԞ���	yx1cSΤs�^?�M� N�cҾR�%��&�bh�!��|+�W%o��Ċ�A�B���`"\��;#��g��_`0���Y��:JJWؒ_z3���J�b�9+�}몭\s��44q�<�<����9`�f��d��������h�꓁z_3����q ��A� `��-�x�NZ� ���sH�<���C�=���A��tc��M��ֱ�������Aϖ���Ť�]�jЂ�<cT\lo���勦��(�{���vv�Q��,߾��+ѵ}|y�(,��̌��g��=p����p,t �O����dv�k�r�Så��{���ϔөx��3��$��80�.�]c�
�IU���\�� �wrЦ2o \��ݳ�h�۱<�U��_�.CU{�tN�eTu�}kwwiv�>��=�6�}CB������!�w���O���_gP���$�V�9v��iy��g% �����Y��Q�MNղ�Sh�ƽ=)���;Pj�����#�n��ɴ��e�'�=�'j�����iVV��s�O9H%Sӭ�G�
zN�2E�a͍��n�n/,����BN§`�j�v�:R�P��q�^`�cBޮxH�JJz6�`�����U��k}QA~D^[%(���Ţ�QNCe-)�e��,������)3Z�4A���)�����ހ�Q9V�:W��"�}��zj�>�6G��;X3ť���W����)�ݣ�r�"��C� z����>��L�nIC"��r��du�{�H]��+>�M1v|�sL�W�4�z;]��:?���Y\F�z��ߩ��Q�o�x�{ҵ��"9�����'B>`����H� �/7D��丼��$pGHf����k��CZ'/*���s��[�>{r)>�l�u/���c	�~��h�
���<싽�| ��+�48#y��1����H�S��d������9��Vie)�;d��~C|�Io3����KQ�?{&ո���
XwS:��L�<_O6��f�%5��}���e�\ͮO����������t�������������s��iO�M;�M9AQ��m���V<ݟ�+.	~a�b˳��Թ��ͺ��ע~�T�No�p�bzv�	s��?l�9/���Ae�d���\J�����Ks�����'�i�ro 4$d�+8�Ril�6@�6ޜx{�Kct��JQ2]"vۥI��罗'ʡ�JJz����C@os|u���G2�c��� O�V�8�(��O��,�?��������i�8��&��RP�z�r�|���N�좲�Z�����I��w�[���2���������MrO����n�u�i6}��Q:7��)�Rf�$�(�������f��B����@�?n�A̩�h$�՝u��� ��D�?G{���7c�^0�t9�{Pf�$����(ɱ�ߣ`}G��}A#���NU{}��ma���;W�6����&j�O:��t��">#�^$才�Ç����� �����U���{K���-Bv�^�++�쑄�����G2��d����������x����]�z��y��|����z�^��~�n�z��|�&�n�	3t���1�5X
F��:�ʊU��Z]w㤉��ׁ7:8�A�l��Ħ)s���B|= *���(S�)5L��K�{�j.�ӏ������Y>3�s���؛JcE-����~Qo3wy���@`4�8w�V�n��ߵ�ˠ)�7�����)�-��,��7���УZ�0�P��]fH�Z��ĤOGB�㍍����Juuu@�H������^���?����1�:����������{�P l���C��21���mDZ4�R2�c�T_���r'U:w���|nre��r�*Z�O��:N�Q��.�R\�R*��"�á����l"��?ɾѴkl�{xE?>YN�̌̑,Hs�1��Y�W��uz�6���I̿C�wR�:"��h���v�.�Y�`��Ĥ�l�- S�( �x3�g~�L�#��:�����Z8c�b����'�C�����%�p� �TEm���~�O��X
��@
 �ڥ��4L�-y����g R�t��K`�9`�%ec�E��\�gh���sd�]� ��V��ɯ����.X� ��9�����]=��5D�>����t]���߱��.����|�-�睹����MMW��j'bq�s��Vō=$�H���2���=�.���s=�<H�wmep��������eD2DB��� ��,�h�/��/���|��f8L ��i?����sp(G���+d���E�����
���D�>o��������#�/�p��P�o�0?⣩���e�����ѝ�w��Kγ]3���hXb��뗙�Tʿ��XY�nk��@�NG�+)MA��fhFWhjd��"^��T���ى�i���@'H>��L-�Ő�{$,(�����Y�k��+(��������9Z>}zeii���
:	�A�������!pQ11@�y���vx]U�NI�.�w�ir̇��tO�n�hVd����҈T��֥����ۇ�[��q֓_Cer�2�8ȗ���J:��t***�?�5)���A�%�s���γ�h5�11�6����2�p��g� �ˠ����a��틍-1Ƌ�-��U]���D�n`�y�2��e���q�I�����������e͑)�H�ȆD(��َh�Y¶����Z�^�׋p�Ċr`T��_&LuV<�./���sJ��1E�����D��(��`�s�amړE�,4L�8S�8���r����#��@Ɖ,L��̸?��n� �����IZ�?;H����t��N�#*�N�>��\ %���aEjP��ѷ�m;��R~2J[��V(a��jE�6���L��3ۊN�À��],E�]�T?���?���z�M��t���Uw���j����ը����Ǉ:>���f���=V��5:Jm+�-B׊���/��)o���E��郗%�T��t
\�� $�z�#*��s����bO���u㖇��6��_3�r̦VaajC��"V|����q�	uuw��,r��31=�K�\k��H�s&7���	����EsQ����0���N	:��
�.H�r�X�께p��UņO��y��~��j� ��T�FJ�������X�k�[���Wę�ݼ/��������oO�Ggq��8�L��1��s�����Z��>C������0��[����i�������HA@�R���?�`��Բ��/ǆ���H1 �Y}_}o���(��G	JK���dJ�@�0�����C>��>0,����VP`����'7����n�<G�"x�7u�ʣ�.y`��|p/�����S� &��vw8�OGsdg��
vyXuC�K96m�ޅ{%(}4�;V���9 H���)�#�@Pҡ|���P��������{h셜TF���9���/����{�1�Dl�g>O��v��>'�}޳`�H)�{K�`@��Sr@8_�۷o�B���A譭�wX/񫫠3 ���O���X?���gO/�_��G��.c0U�!�:�=��tm��S�y�<g���3��\��@:�&*hiYH-y�"��뜡����K2�;O�	5���!|24� G�邎�,x��0e�����������]��܈9�OI�Y�_{<=b2[�z�}. 	�'Ř(�y�����@�2&Vf��F?w"��g}��#Ihxy�7Q���U���|����z��]��V���;�#-}������y
�����ҝ����/��(��Y��j�@�ͳC�&�].M��EеB
wSJ�,�ISFF^i*0?T`�ghs����t���pqO�0��!k��o�j�X�8��|�����Wn �l����C���F����'�9L�=>�À�y5��~�%Z���j��rmn��?�9u�T飒����d�>(~55QA23���f�eq�f����c�HY���[�]���o`�cx�[�������x�sV����:�Toan����^���(D��	kc��I�+�i�
:���e��S}��a�߾���Qκ�du�r$bS�w�CUaӽ�^��j ��o�;�&s�ҦL�E��\n]'������k;�&��mqqq��|�f���Κ�׮�KI9��8I�'�Y�?<�h�:����*����W ��mYY�!oj�� ?+�ٷ���)S4ظ���e@@�YR��@:r��1� qdnsI����%G-�����TW�vxz�*N�H���2!/��e�C9*��n�̨���\��o_��dk��L���)���ze+�ƭ���Έm��s������?�����(���L��O�?~�n�	{�
et �Q6���޴��9/���'���B��A��y�noo���B��LrJ;�@��!�����؆�M�����	�{6����D��G
�Ϸ����J�k'�sMinj
��/�Л+)�N\l���!�"����<���!7)fcCX����,@����S��1%7~��↳G(X�_��U���f[���²�.8b�Y���@.i�\[4܀=������2){��>&��Z��EEٮ9��s���p��s��n�a��-�dR��ӿ����gv�˟��E���Y$��r�L���|}�**�D���7&4�u��^��Qʊs�����6���_�;��.i�\�$�ɕ�_��NOO�9a��@���M	ـqS�h���V�89��H�W��=������u�J[�/��G��Xn�?Y��g�X���_�[xV)�}@􆷵�!|������!�:l�6(=�Ur�O=�x�N(+�@}
�6N�am���3Y%=K�s�熬J�f������F(C��Kե�L5`���Y�V�=!w�	�����ɻQ��_��?�Q0y�����4�W�ݸ�z�\k�Kd7�E�wnu���8�{e)�#KJn�]),����;B���:��s�HQN1*丢�b��*Љ�/��&�&m��7�"'�j����!�b��߁�����w�o�鲇ؕ�%K�bOU�ggy �1�=rx^�Z	���f+������.�-�"���m��w��BC[��=E

0k�캟����}�����,8j��-l0�G��5��Y��h�	��)-�P���bL�ܹ��w���bw������"G��1�8=�����)�Db��{��
(�ܘ��g�2��+qW��h���� ^�ҒΛޅ"Y��$��Ç�iԽ�ː���TR�%WWW��Z���Z�FG_� Q�,�!\�9��OZ�x���Z��v4.���f�y5z����{d>Ϲz�%�X�Cك�kq#)q�!gu�m	B:p�l���x���4P��-�ꅚ=%�xע���OꌡD@�#E	�Qv�O��������x��.����l���ɉ��f~��D3���P�j똚�jk�l�*9y�b��<oj��Ѓ���Ҭ�g)S���! �0�}�h&�����F|�O��z~���<��sl[KGx���5F��Up�+�5�7o��¨U��Ռ���@]X�<5/`�8)r<�7�B��|��.��'�:?Y�}�u:�%;�� ���@��O�~�6�K�!��J�i�D*7��t��uZ��˅
?�'�}�ś	TT�l\Vpێ�2L�	�7�4ܜ��n���;���ə�z��I1�4���H<h��4�XQ�xQ&�W�T�����KP�G������ӱ�F�}ij�E/l?�XU���$
�LYF~4+9"�m����ש�C���a'��0���0�e,��R�@�4�`)@ɾ�E�d���'9�|�h0��������øn��:P�����5���%;/�oM=ܽ�\��^�Z���	ʼ��pq�2�{�;?o������d-䟋B����%qiX-&�D�; �͓C��=�$��xr�}^j�5&ff�-�^?�����)��Y��r�T|P�Ql��O�K�(�ݿ��'��Н�V6�μB<�n���W"r���=VA�yC/x��W���a���9/�)+k����oғ��	j�
y�	���Ŷ��^L��(��`���o��6��rx#-Sje;�(���/4�6���\������I�tOL����HJ>il���D��AN��QEy�\\\�R����:���C@ְ3��U�1�8�3���&U#��S"�]��<ćG�Ľͺ�Q[88�B�s�ѱ���j+v�{g	2���m�uHȥ<�o��{{�Z�e��I�$ht~�wA�]��z"m>u���1�$�rݸ�����Ѕ�̡�;ZP<L̄������f㈿������_Q9�x叕��]�h	��Э #����o��gM�>��S�#-}�8���:�{su�P�К��ܸ�Ljo��8*Zu֫��g��1RN�yv�|�ghx�B�^oz�w�{2���i��%s����*=�����\���c��<(a �A�!��=��/���x�0yP���fi�(#S,R~)�	����{��A�c{9���xP�/xe%���A6���>f���%~��I�U�K+��M�J:�!�I�����z�LHXCO�/Z�9�V}%Y����������}y�.�cඉ��oK��G;w9��y�fd����\LA�k%ā|!**��4:kx�̄;EE�A�ϷI�#�Y�� �i	}_�v#VTx����g��HZ`�@���G����J��ϟa�9 �̮a��z�����W������h��M~*�S=/��	5�<y�2Ug�N�,�C��vB�5���w��(��*�U0|�pʯ������w�
>�ss����N-���hW��[{�sp|�����6@�d�tKg��E{��Ւ#^���<�m������{�A;;_QU��4�$ޜ����aw�:&��z�êo��$*�E���_��L�����HP���&�!ߑ!��Z�*��aO\�ґe��k�"��'�G��\~���^���G#yR�x�ī�3�8��S�Hz��R�a��Bj�H�O��E��~�T�K�Ջ���>h I���B����9�w(��x��'������E�؝�
���:)t���	�s���D�+?��f��IJ��cl��V�� �^\ģ��V���ua�����_T=�
��l�Ƌ���0�|.ךxv&�Ńx���r����t���P'����&t�8�������'� ��)q_���KA�'��	�̄���D��P&��1�����Y.01�$� ����X�T��@�OZ���@�ƂB^��	��B�99n�Ԏ�2��hDs��A5����,,����~w���-$�� �蠂�w��K��.x��?����=E��wx8��TTJ�xW@R���5�l[KT��ݦº�����F^��Ew"�oP����^T��L���?;���/��q�ܛ����B^&W�T�IO!�uś�%��4z~R�@��
��l���Y����<VHA�u���_�{��YJ\v��EɦS��TgζbW���:Y����*j�`�����nH�R��Ֆ߸K�ᠽ(ݧ�����Hԩ�m�{t$��m��������I�-�?wvh�%|2���Q'�ez����	��4�d�֯��p	0.P[�c�XR��Pyue,Ql�vC3Eo_JhB�j*�{���s&��G�O�~9��w�`6��UVH��a��<w���G>F����:E���Vx���FY�03��R�֖p�^���b������)7�nF���G�k���#��#�e:;7A�0��n�ʌ�+�������K�Mh������6KJ�&W��Ս��@�R}�̮ޘ�|��8[��m�QW�;��/�7P�j�R��1�-���t���'�7,ͷ��PlZ�Џ)r��~�>ˊ.����/2ά�M	7ZA�+W�\�E����=��0ZͮRSR��R։"F�JbM��.\�"q���4�s=we�z�&�����q�řĦ��y~���aG�*��8h��٩�oG#c��7u��?�(}����f�ۺ''� �$U�v��&����yNr{D�!NN?ad�?�Q��CT��������φ<w[[�n/h��@]t�7W������[^�T&���1C�t(�t��n��w�束�N�p=���d�4��iK�Á�����Ev��]@�鹽nA�gٚ�GLb�6�4[��9��&~��u}��p%^-�����N�q	�X����`e�V#������o���W`��ga�����[��geq���<4��\d��	Vnn���6��wh�`�`�y�� ��*����B��,=��,�r4���r���b����s��>��XҋI�Ƨ��G�� ��x#��9մ��+��h�N,DCHo�wB�n���4�-���������=yش��qh�;d�o$I���c�x��t�dE����j���E�:��TA��^ ��+���-O by�RI:F���a�Z�|�:�;�4����)ǯ�z�����p�q����PQE61�6y5�b0������Ǹ�:낤�ʭ�,\�8����Q'!�8�K�l�
h>��N��F��8��vu�<�quv������.G���Ø]��Գ�'
G�Eu ���DD'�o�>:�y|�ʚ�g_]S�����Vi���VWwwMuuDM͝o��5��fA�T�뤯�()��/н9��C��y2�G�����h�D�p�e�?0+�H��dH� ��q���P��0����G󾚽���wY�x/�s��Wز�ڗ���;�^���m�Y *o_>`��>����0�Ɨ���汍&���i�ts�����<�
����\t��*{>鵴�G�Y"���������z�k�>� ��8ƫ~�q��x�B�U�:��[�K��"{��MZfO��w�݋<<�
��Q��Qо��uLO���c�Ѫ@�;���s�I���+2��ױ``!��(�/4�8�R .֦�x�$�����b���̜��P���Vl����i�j[*������EZ�55
�H���r��^�ٻ��载A�T�Y��Q�zE3�m����!�3��o"���2��2@C�@R�K?��B�� r�_�;�����H;;j�ܭOn�:�_���!�G::��\_�20�ii�Q����b����`z�ID��&��g�	^��\4�ZOC�wG&�$O�5 ����� ��$B��a���m"hl�r�jn��T�����?� p��ws�AyGG6�Jd8U�x�Q�|q����XQ1�1*Yl����s�.p[�����Z�8�`x�ocZ��J�f�f�}���h:65�e(�	}���Tͺ�N��=��e�R����bȚ�~�i����Qi��ʗ��
�����+�́%��d]óm@"����H���rw���Iq	�2Y+��K��
EYRF��{5~�^�+��{�s���j�x���;��"�bG�X\%���%g�Z���h�za;�>������+����F�
]2Ck��OשB�����d�၀шB�8�!0,��B}�]����.������ʇ�C[^��[�_��(���ߖ9�*�-EC��Q++�H��<'�WQ�*%����
t��(�?�:	�*:9�`u"s�\K"�kqQ�1��9���}�]��ZKׂ��d��ß�y�������먃o�_Zg*]P V�v�gz�u�<���w���yh���2a�G��<Y}���lt��Z�x�~��*�>̇A����:�{l�AJ���61��{l�?x{��$�Fz�U@����ʧ$��۬eͫ1���4,Nva׆ �v�5h;=&��tИY[�c�t��@݊���T��ɓ,J^k_\P&��Z��׬���q?�&���%���?�#%��	͝L֣Ňn����\wuo�5�E]U"���ż9��LIDe�>���~�)M2Whk��%@X� ye���;Z!��N(�2�\�����p�{#�%�0WUt�̌Q)�B�dk�X���[�Fme�H�����A:��?��J�q��� $Oͯa3��l��ͽ~N��������Vw�t�1�r~)�����b�N|��cc�Z..�:��4x�0��蹎�<��uV�aa�noϟ��QR�����ܼ�%� }TZZϵ	$:�P� �9	 D�R���0���v����~���knS;��b��]|�������1a�d7��Cc|��R4Ԃ����G��򱧨e�y%0��d���bç�m
�-��������&z7K c�4b���3�H*8ӡ��r����Q7�+W�FTW� S���q�/n�|2����,��������q� �yFF�ی�q�y�z���.�Жu��#�����/��<��V̝��<�>��)�@��0Q%�0%�{��i��w���I��aj�g؇��̢�f���v�:�ƴ��;'�Ko-��.��/e�#'3���TC�
�\���Z>���1*��c��9�?�
�Nf/N|�2��Z�x��tR$v�'��EM�.-�9��Ң\7��CŁ��b�!A"@��KM�������?y2���j��]f!���DD����X4��a�J%W&��G@�1r!N�2;
LU�.z��v��OX��2�j�+��jddb�Ax�[ª�|}W7�TX��Q��Jx���E��x@�a��7�[l�M@�k���1	-x���Qҏ�^A��g� ���[��4u	>9U�?��oX�o�x����Q9��4u^6����	\����9��PK�,s��8��B3�]��Һ�e��Y�0ց�TnS�"�ؔ������q|-���'�/J���6]�&@��[$�sf�	JЌ@F��]��� L������akg�R*4�5���	�#�Y ^ �D��tg��)q�"P�����u�q/��u`�yp�g�����`�+���ˏ`Dި_�L�����P��慙Y�c���%P�#5Q���Dًh������h���Λs~�_GA2R����p]�OrC͞��tdk������ݦ�\Dkjj�����1�VϞ5V�<y�����L��-M�LbjjS���h����cq�� H. !T5���ڄ5@	���|=��M��� eحS/KI���e|?����t��WG>Ua�z$Q��Lͫ����&�Zf� ���F*�S�J�ms�oǈ�k3FB=����U��0 ĺ�~�Wq����>G���d(�����>%x~�>�	�L�&Y�
�� Y�#5��0tJ�/���._B"�����QR�5��}��vu6��i�g�-���'4�"��dXnecCr(Z���#��6?�U�	�b���`����^��i�S�$��NQ�M<�BS{b���t���?.����,�٫"��\�7�p��	rl�5�I��_�H� u���{��T > gi�l\_�܀<V�� �i@�h@�h~��P�Λ�� 6/f�%�%��6�w��VD_#c�
8�NM�,h�s	bN�t�-Q==7� j��;]J�ƢY$�����T���,���u]�a�� d޹��nm;U�=1!�G�����0H�gte��Md�,)9).-=���b�rH:U�ݺ��_��>{EaEA:�f��glf&��X��ơn���^�!a������y4IGŻ��+]�/>a���[=���/ŏ�b!���B�ZOL�Q|%���*��CHJ0_�J�h�w�UQ�2E�XBF��9�ZN:o���h���ޅ�߿��HV�k�OM�y���}42k&�F��ٔ귃2P�DB �Ld��˄�In�J4@�ҦU�^625���P��<(+������6� �b-�<|}���s_7��IZ����,?��c���^P����^��TvX۔�/�o�o��_���>~�B�`rn��N��h�6���� �#�w�U�Q����' h.�U�5*:Xri�� ãY=��N	Y^�(��#R� Y�Ȉq}�*� WXH��,�� l���&
�a "f��`��� ��z��`3���o߾Ex�֕M ��������_��q%�yO<y��Բ�] 2@��j�����a++��s�Y����m@y9ڊ�
tD����sZ�a9uH(H��Ľ��OzEi�y�h�b�c�Z!��u�j��}&�Ӡ�uD��Ec*1�'�E�Y�"fXo��r��R��ffe9;����_
��EsF��0c0���k�W�Z�@F]P SSS
�"p��j�7PPL,�Q��$�@>�yKH$�I�u����7�t7����￢���X�B�$���>{�_ݣ��C"����P��Y�#��J�Tu*B��i� %�1n��=Rj�'�@��5![c���|.���E�V�Qˋv��5_U��Q�\�ʚ[�5���;� �a�r��!�8"�1"��CE�DGWyz{�*p >.�����14k�I��~�%���#�;��������mݸ���&�@���1�VUu�&�]D{o�B������}vv�m�)f�^�\܍�zg4��a�e�|���b��������ݥ�*9��s�Aa��!*��z�
�J����`7o*x���yW�-� �K�hBh(�m�{es �#�{�~�P#��:K(r�3�E�
QE��B�U
�0<J;�������3�=W�{p��]�����Fr���K**H����ﴶ122
���G�A����Xb��5ו�ݮ��5wZj��[[��P�;HIE���� 8OVO*��à�����q.2E��ꌅ|p��>�jS�Y��3dv�\�3y$�%/�p���-P�~Q[)�z��ǘ�& 5��ԯw�n4���7��.��2��\�D�ݯik�{f~g�A���M�AC�$����Y>{��qٽ��f��v��-�v)G��{�������M�G8[[S��g�O�24,SZzG�u>���b��7EԜ^`!�:..�5Ů���-d�R�Qb�u�4b*+t����a���@:(Q��A�1��)b�/{?����¸N뚒�m-6�\������a�	��Ɔ��g|>~bwx]�]J����K�NDq�u�\Hb�x��\jG�� ��X_X~��X�߮c�J��`#*����n��h�WJ����d+Ɋ�N:0
�x�b "%�졻���T�7C~/�)ll4�Ѕ��s�ܙ)rd�z���"0X��|��Q4�~1
@�wAӨxZ.��< ��� ?�Wq����+$s!�@��{��l.���U䢸�$�����d�a�H�I4�l ���U_I}���%a/%�d �������xibn��t��g���=�Z������l��[�Aosr��n/�nA�p���u{�y�����-�э�h���\��5��B����/�y����4�{��&��V�9>�$-�8	p�� X�Y�{C�z�.5!@!OBd�/P0$���:�������'���b�}A�l4���4���v�`H�{��9�7[� ��T�� 1Y��rfX�D��8�9�o� ������1�R�(+;zo�7մ#��'�d����Ҡ�y7����ܺե9DHS�d���b.���&?+�$�sJ�;�g�
����jj�hCZZ*���ڀB��H\  ��\��?�=����z��z��b2 c��k�'�]E�C����dH��� �ygY3�0œ�v���hp �ᢈ���e���g�.��+�CENy����e�LJ۠�*�|��ue������!�)��Z3�і�>أ/���8)�˂7߾�W����8\X-+�,8�
�����X`��/6�T�SҎ�x⌌�#']Q�X�.ba���?���0�ǻ�&��3O����
��)U��SJ��ӝܮ<w��ڢޱԑGB�(Y�h<T�<$̪�]��oc='���䩔��~��6�",����H�{)O?��=�'��+�ͬ�Vl���u&@̓�-.^H��xp�?��B0�Z2[���ʛؕ������c�8R7�A�]�I2�J.��
'�G�T�YԎ%���'�hs�q���32"�
���;�5?Y��"��Ġ�T�d����{|; ���]�L=(��7�/���7�L�t��i�NO��7(;z�Cf�y��s Aк���L�t"f6TA�����2�E*����i7T<ծBa7�:���hq��龶��ћW��؆�nˌ8�wD��߄O�;ՇyeT(	Kx������k����_�8��Do��M��������Wb��?����;�vS�R6M�(,�C.�kp'��?�.�ך5���[+���֣#aqf�9�z�M*\!'77�,���S�-&�K�C����d���OH�6���>��b^����zǦFq����C��_��R�s��f�A2��+T�d����| ��dfib�����l��D@�dr�,���]�Z��W�9Z5����Gr?m�t���P�A��{e�Nkr���Zh����o�H<*���_�Aߘ�l�*���A  X����|�'��u����}D;�Ho��j��]��<�r[<�@MKK�M�/W�>/� �3���_��6]����g��D4(�����A�(�J=i�a���^�?e���,�a���~MS8σd��������Ө7��'("PS�ޡ'�q_A��p�,w�����<���]V 	!i����A����5��X�4ܠ��o��%�РC��ڪK�>o��	jb�;����M�ȺQ&W�&�����m�K�擗�����bT$��q++�?���^~A_�D�����}A��2�Vv��U6L�!�9g�Z�|9YX��yR��z��ˇ�::b�d�_.���iॿ��p�<�H���{�w��S@�:���.+�v;M,�~�\Nظ�0�s$��!��UN���&��u}�E�=�8HRM�U��B4�!w �uFrR2����o�G e_X��=!��6�V��Z��{�H)+��rzZ�իi��?�Ԉ����q%\�%�]$edځL� �[B�A����p�d��������r�{�Nf���e�.I��hL����G�I(��j���>���1�MBA�_̄����F�T]���bE1Ȥ�q��>gı�ˈ�7\+ڨO���@��[R�_�z�r<�w�sUmN���Ag��|^�:- ���d��B7�>O�?UI��X9��;�Ź�t������
:1y�[Vf�=�/��q�n�r,ad�+�����Z�������$�m���D{���Y�˷�_C[�|6.|� �d��޼�K�	�&n[cK����3.(�
h?`9�t.P��*Ε<�,��x�`ÿ|��,�^y��P5�GN���s�Ms�����A�7ڡ�OZի�p/e���)�a2c>��3V���j\�:q!H�:E�埰V8-�� � ��z���'��d��E]uu�}��Z�~��h:t�Y��Xbjj�Q��e�33w٩}�y��b[�˿��<}z�P�,+ͩ�]%�C�k�76����zl�V��:��� �����ꇦ��Ŧ߶�=8����j�A��Ukv��
ex�)�<���]��n,U���
i�@V�Fӆ�sv%c�{���,E�|H�x6��)�l����( ��!�#�ҟ���D��n��>�<a�v���7�Q����w���2�;h#=�[�?�-��h�*�K�������T�7���\�Z}}}�L���6����1�6�KGǫy�%G^�/ww�A�C��[�gϨ�,K���쏏�x��!Si�[�q���E��oH3����X
Fh��j�A�k��є��~{Mc,�<�<AE�|ԟT���/7�l�'��i�d6���n�]�Do5M��L���?�ȉQ�y���wx�|d�}�Hd�\�]�� �ey����*��y^Z��4��b��]�%�e��Q)����aL���{�SY?�5�B2+9���w���}�إ2u��Ʊ��V�=�����z��Ւ_��6m��.m�sq������l@楥� U�Y*�WW�/. ��W)�5p�鱥�mBV�۝���d�F����.3T�׽�IE�(������7��|��D"GE�.����xɫ�Wc�ZO�Y��%@;H��̀����R;Q������Ap�
�&&7@u>8��`e�G���쨏4��pZx��Z��e������P R-�ˏa=��RL��kC�`�Gp��b��R|������̏3��-+�(f��VV�=��11�V;�
mڥ�NA7�B���8(1`�@�-7���jRl~�F�&_�R����R`'�O��vE��	�AL�E5����� � �F\��(M��q��7A���f�`��DL?a���]���r���Ce��ޅ����؞��饋��,��g�8�_ �_�я:-�����[�>�4�ǀ�%<{aw����e���Mc�2 � �t�����_�ܹ���zw?�;�;���T�k�QiDx��+޿ק����ո�|��L쐀W���-��b�����gg2�_��
��u!U�z�7���hv�~��q�O����+�~V=Qs*+.�:R�R��t�������CP�+�/埇�;��g]c�+�l3�-��6�w,�Ot�.�$P�77J�Mp��YT`Ra���!SԾn�졁��0�t�\��g��\�Lߵ�*���g�hb�l���x��j�!������ޞoU0?7�2NS]y-َ�oc:����d��������gR,��9�-lm����_�n��w�1p���	1��Y47Z��sjj��P3�֨���VKojf���_��1��[ʠ�a#���,�J�!�Z�X�꣊!���"��Gʈ��S��e�7����*���KM�����b�kh�����i�/3%eJ���>��ۀ���{Ǖ�шh7��� ��M��8�L�Ԕu��<'j���}���L�G��D���ٶ����/��?��O>��W^]_�=U�R�]պ �v&.����W��������bm��=� H	�i)�s�0"���~�=��^�2vqu�HU�ՁFuZ���{�i>��_^�p�a������-�5�T%*��5_$�|��[��px��[gj��k�`���!*3޼�H����2��тJPE �3޾�9J�r��˂��0/(�<%�ϛC�
p~���^6���:�\�L�eM9l�n��H����>A{+7����QT��F��l\�����h�h kfN�*���^��?''E����y"
����Lk�V��~	9-�4:�3�B$�h� ��Iz3C�;q`���
@��}�l���C��b`)�'Εչ^=���2y�.��v@�7�B���*%���D"�k����EN��n���^h <y�U�X�Q�ܢ�Dux�44T�N�6�,�Kf�eB�pA ���yՆ?9���p�0F�"�pf�;�
:w��\����UX�,Z��2��x�d���|] ���?;y��{?@hC�)⿺$�%���C��ޮ��O
Q9ߓ��͔���Q~��dw�-!)a���:h )촮�X�	=>�� B�Y_��]78c�O����Ԥ�Lv�"~��͸ny�#�\�ɔ_�is��oQ��^R�%�+���/����GT��/� �ɇ��P%g}!7��A�`�V�K��N�P*^��O�i)/CL�-$�FM�ݹ5<8�Ü���n@U,AJVS[{��-��J���
�D�9�}�v�vǁ0�Q�H��5)��\_'� p�\J0��=Ϭ)q(��
�{�@�$@ہ�8)���d�	�����9P8%e�F�59��w�G!�����������v�|ȇ9C���� w�FS!R��1
������tt�*�����옟o~��Xˇ�Hˊ�n3)���)v���d���vw4	wv�Ǭe�K���z�162̿���ՙw�q�P(h���̮.�������@v��k��cuc)�^���<9�~L�o �(�P�'����؋R��X0[��5A���\�����2Kо�L٨����6O�5W�%r��Q��w�A�e<�rswV��ꋲ|����b` ���y�t��i��G2��R2����\��E��<�:���1�>�L�j�x>�x���s��sCFN� �}�q��G@6�5�����	{�u熄�S�v����VW�X�m�{2 �`mk�T2k�f�F�+��"B}ȁx{��UÃ�Cd��� dq�Z��/q��:�q�A�S���t�޸B Τ��s"�29�:!-d�
,}�u�7Ksuo��̙f�����0��S#/������'��H���
���xi��	d�z��X[�0t���<���12�����1D����M(��6p �Qm
������&S��e��a�yXN`����s��&AJ����L���Vf��W#�cВ���|i)hkt������Nn˟�o�G~N/d���9=O���Z��^�\ĘY�W��t�r ^��W�A��/:9�:���\P�}�D���m@�Y$o ␉��7s�c��� d	j�&U�O������,�Y�C>�]� �?��RSS��=qIX�犘��5᳏��g�C����ie,0/S��-�w�0�F�EC���О�o��o�UO�&�;)t�6���.�΢,.�sm�73�O�ې��'#��M��1��sUv�gb���@��;�����zpy7���ȫ��6h�1;!zPR鴂�΄dBH�����&���	-��K�V��_J[�Q�d�E�o���(��-�5A-�->�5!kO{�Z���/4���/t��d�ok�,h?��������Vܿ�p��J�^�zk�E��[[��������>D.
�fFF��!/��*Y��ch�Z���GI@���|3a��ܜS�il����>��g������&���hY��>)������34N;�U)�:�V��v[>�ܾ�HK߀�iS�7�-{X�iH����\�@�8K��ѡ��7)��Ҁ	�}7AN]���b������V�F�K���Ž{�z:-�����X[_�1���kfF�PwEK��/��U�8[��OQP >ǚEq��H�ԅ�9��I���X
}���D��d>" �1J�m�0��@���;������uR2�6���Ҕ}[�йq�g��29td�@�����9D��nSn���1�<�Y;%�(�n�	�b��;�q����̜N�g�eN���!`X�R����ѳ2����ii/��V��5�C��y�՛_)���H|�v�ʠ(��f�*�ץ]�E��w�h�0	�<$2U,h[��Y�=���,+�=zKԕ|�V|�妩��=��ɵ=��n��+*�*4�9�̄��o�Ǎ�ߑ�&���i�+��v�}�]��Ɔ睕���nϥ~�OO�����3̄�Q�\}w<����$Tv������QfF���{d&3�C:!������qp̬����~�����qz���z]�s��uߗA*Î_S�2�͝V)��s :G���	Co; ��x���ڸ�� �ǫ�w��y�H'�N�-E�с�#�-�*K�z�=�sʞ���s��N����"X��MOs��U��%YA�
����-��?�9�@׏b섳�:��!��Y�h��{��.V)U���>��T��˭����B�J�	�^���E�_�V�e|�W��=�����G; ��'-䵯�r����.!�3k�r��������Y�vt̼��R��y������/��,vq�{�sT�_CDY�a���è���HVF�����DD� e&`(Pd4$���n``�^W�����Xoq)�*���,+G��wO�D 
Ϝ�FZ+20 ��|h�CS{�G��%��?��|��P�H`��v07�����e�`��y�q�z���<* x|-j'����<��aWWW`�0�78s\*G]%�\�3]%ze~�T�ԉ�f��5��WG�W�z4�.�w7cZA�����c<�Mp��b���9��U(��N�b���������,���/2����?���"�l,�O �L��C ��(��T5&�z��$01����$��Lֹ�(��z:���>�����O��+&;^���'t�d�hbPӗ�6G
�d����H�E���N~�%�<���K����ڳF�s������݅_�A� �E�3�c٢�ed�����[ncS .�ۡH�`�F��D�yD��,X���@�����Ig��=�@�d��߆,�ѯ
4l��6�0v�G��:�ׯ%�uӳ�Z��ǿ�ml�����=��4+���4Ӡ_�r.�{ֹ.�r,��Q�Mi���D���8�VO`�������d)��JM�;��ݯ�W����h|��<3��o�Wֽ���a� �1E�ܼN9\N��0=6�(�����WE/4��]/�]	���f��Oc����p*�.Kʚ�Z��;J)f�>5�jl5|��s��p�mb�sJ@�s��yO(��/�qwR~"O��ʵ��t���I0[�����N�M��B�EDkɩp����j��;lji�
j��z��eceDZ�ԭ�Z6�$�t�{�\�Mu�Wl�^�{x���p#�cq��JI'�������A�2�<Ԣ�$��nݐ>ZIʘ���]n���k�*���ª+��S��CC�f���M���߽k������������#�1`��w�F|-9d)��k�kR��~ڻ�]Ž,w����F�S��C��q������Q�S5��� �k�'�e��hnȾ�a�"��E���'�o�k�����=�sR�a�Z�ǥ���b�g  ���mY��͡� ]��s����p=�O��+��C##�h�FJ4�N�s�K��'���:�4�u�me�DV�7�Ȕ�0�C����@	�������֒�Q5O!ͭ�?,K�n�9e:(�jE)��D�nLq�g�J���q�m��|�|�/����S���/�#a��;W1<:j9;�hE5}>s�>u��oJ��Hx�M�%	��Y
�]_�VY��ATy��8d�]���ZT���sV*���c����\��(�y��y�!x5�;��<�_�+&0HeW��y\vF[
�'^�&Y���ϫgߌ�O�'�Ϗ�U������Ĵ��F
]�W3�Ǥut�b��)_�'@�U��:�4퀽����Z�D�$9t�HʣK@����5�rNE����-7��.jj�VnF?W��2^�����Y��2�v���c�r��e���~:�\�6.��NA���|��٘;��c\�Z�z��AHh��7r���tj�Y�s�.��:�/��#�n���Z�� ���V����=&2_)P��뷉�!��C¤ �b������}'�Jy~�����*?�VTN:n�>���C��8~�%C�)����(oK,�������G
;�F�����%%J�����D���R z���R������-5E@�;H�+FHD���GG�a*-}6����a�`����P3Ƕ����UT�Dw��_�φ�$��x�p��,��x�Ĕ���vg��;/>��`۠��>��Q��\ZUh���w=;�غP��Cj)����w�����i�_��/��!��b�̒\u*�w,ohh��G��am�<3Z��̌u�<>���W(�jf���%*�!z���������+�^�O�&e����O����h���}R�k��QB���+ޒ+ޝ�������GHG�e��c�m/Q�� �^��ݽ(��%�g�ߙ��K��F��t��i����J�Zb��ƀ�^����j 9s�DJ'S���[�Ul�����;Z�ij@��rБ��7�
��������yyfQ�� d.)����s�����ܰ��u('�����9�r� ��D�=M��wW�ր�C���N���@P����`�������e	��C@&-���F���"���^TD�e�)�_g�'�F�9�ח�|����؃W��i�P������#���]^''d�̢�Z�^����]ԟ�an�OPR�� Ds�������ŏ�O
�O}�1P��j��E�;8\[���^{��iG$\C��/5a<�-˻�J��\ިQE1�{�1�����FC�� �fB��?�Rm��~��U��_�wׂ4<�,-8�Qt2KP[�ݻ���Ǜ�y-��j֮�7D��B�Ot��į��D#jk�Uy���E$'�=T����\�zqZ\����j/+Z?A��<k�n�p�9kr��8��ߝ@�Jw���R�ՌM{JL{�M��O���v����J'����is�\��������ݪ�rrbl)T�����;��=�<�ۨ�q�).k| ~����(!��E��=�����Ef�뛘���/7h��}A"��եb���j��'X�(D�:~-2��o��[v����"q�ؙ)�r��I.#��{}}���O��3^���B�~ �KV�&���V�y�0�upw�F � ��+�N�����]^����7#�`JE5�� ��W�KV��\l"^�Aj���r�ו2���b���z�� `�̤M/r���pE�4�j�U/����>a]���6[f:;��ͤ����KM��o���hxX��������2����9Y�;:����T���=;t{��S�����:��9�ǥ������G��\�] ���I~֭hJ�H)s؃ؙn�ݨD�}P�{�)c��ta������l�ݳ���;��{�AK��Nv�41͘��ഇ�<�>�C̈́�%��Tڝ��]<Ƿ9�6���SL�Mm��e<�z������f%�h���A�^�^pչ�~��$�����aj%�V� h�8�v^����խ����Р����|�.�8��d='~ [)�a
d&�7ʇ�f67M:%� ��XT�}q<m�?�	r���j�w��Ϗp����Oaj*��e��D�}�e����?����|q�~�	oڕҥ�5�_��; ҳ������,#��A{Hsf'����\#� p�L�߇�S�}^��]���{�S�9�,L����#�HX<)?$;�QJl�K���fJ�(�|��x@�,�.��_���뿥&����o�8I[�$�2�5�,��E"���48���t�����!�k�������N�X5�^=�K�b֑���V�G��_��g��yeO��Hr�:ryO�m��6���Y��j��;��|����g���+W���Fi��v�&�����E풒N�!���\k��gb��&�7�ꂃ/dkڎr�OO7.��$��╦rrp�5G %��O�*Zo�d���=�A�s�@�F{Z�}�T���㈏RR��Ώ��jν;_�R	#��t�����%�/����)�d~��fNN��n����>16��M�<; %f..DYd���=�E�����&�#��K��H+'���{C� Z|4�AA5.�S��O��+y�P���Ž{�)\�f�A�d����U���	4n��BJ��Lx���EeX�7�~PAԊ!�5�}���	(+P!�J���R��f/�fD<)$q���]5,����6'k�����л������G7ڞ���x�]	��XB/��3xI�?��V�O}�=��I�W-¶��ϟ-K�q�aI�e؟W,uu�c��g��ޑè�:�oN�Ţ��d?W�po��''u����ޙ��B���!�s���%h��4NL��%Le�w��� �X
|DP�R�6���+�K����g�o��V���$������s���8��m0)+9C���
3|�:@OX��Q�J�	�y9���ޅ�I�l_J�NB�kb�FAƦ���v�܀��~q���,Fߧg6	��b#F�u�B��BW���wg*{�#��H�(��x�9�!q�dnD��|h�݀��e�mtTDuÉ姽��.�������$���tJ���`����uꚩ�Օ�EZ� �O/��4Nt~3y:��K�e�0�	��̐3,���Y]'������S��L��D���Ү���'�
���YY���i��N�ȿ|�Ni�_�",)�8O�]\Kt[���G �:~��{�<�B�9�(�*W����@��Z�)}����Y�|�gKo H%'��Po�Vґ�J�$j�{Jdm�(è�L�˦�T�><a�9닅U��Q�EF����޽[�����m_Mc���S;�qеpܿ{��w�� F7��Q^�Zw�j�I�ϟ��&s��P�k}O{����`�rT�=y��J��'��`�X"PDiC��FEE�}^��[(ޜ�M�	�$�ɺ\��>��A�Fh3�\�����u�ե��.*����3�/UL�[F���T/�� �U씁Wj�bWW�So�.|�7�Y��x�E\Q���1DǞ�U����ɑ���D�Y�$yt�q��r�)t.Te�Rﳿ>�6)�	�y��2��\����V�.zջ�!¹��_C����G��N�u�zc<�ؚ�:B*#~1�D���u�4��ܛ޸���,y&t�v����H ��Ԋ��Fj��UK��M8/��m��z��P�r�f⇶ ���ڳ	���>V����^�z���Pm�U3[��0�����f�7�û�1�(�jNr��G\�fC�͎ �z	C�?�����dZ~������=3#o�am���vu���� A��ϟ��ǜ���l�9�3���751Qc���h�}Ë������.	f��^�WK�X*�r�Slp2Ĳ��4�җv�k��4.|�U�w0���R�	m�s��E����2M�7�<�^��e�xZ��YW��O���������	�	�Z��:7/��M��R@:���ȫ���0/��s�*� ����\�(W�= ��k3��t-�wW�FD�% v6����M#�\;~)�/MHٜ˂[7�Br ��I�G��bݩ���Γ���X44s�wה�|w�q0]��]h����\Z����:`�7�g��Q�y�<a��:�WVW7;`����5�Y]ݸw��1�?�<�\c�T�i��K[������P�RE嵐�}|�V���F�J�`*đ����XRSSe����B��q�=Gy���߻׌J���"$�^�%c��gT�k�Ɯޢ��S�YY9�db�eS��JTy]W/��
�����ꪗ3ˇ��~GQM>�+�g&������!��	�1�/Qy�B���h��'47�xRl)�NMo��5��U#�m,�� O[׏��_��M*�P�S� ���b�f��'������hs�3�Z"_�[H�H�M{z��JD��e��D����K�0����fA1!Q��4?/J�(X"y��"W�כ����8����w��t��s�WK�Ͷ��p���^ꋫv!t�� J����H̀|���g�3��&O��ʪ^�}e��8謋�(��J��w��2������ �m�[��k4������$�~�@m�Eb��:;�^~�M_��m��]���畒j1 �E/�a"���5�����c{�tLB��#9S�A�����MDX��JKd�θm;H��Ꚍ� ��o���BL��\��ۯ���ѵ
=��х��!'�UJ�n�M��%f��#pK�b	3�źF���$�4��EF����j����L7#��_�+��Y��Y��2C�^�23�zU 	��HB�t*jx|\N��������ȋh�Hmz��lQ���d� 01[e�SS[�u�O�ҩh�S��[X��ݞ�6�7Vw�9XA@�5y��������1@&�����,��S�+���1d��S_��W�#1�\�0�� _��#E:Br���Ն���W�Q[�h�P�\sy�C}������d$��2Ԥ�z%z����5%7���
 ^tRUR�����Գ���J�g�J��G��1��
���ۻ[�O�;N��������MM���KM}������V;~�Ș#�nm�2����	��qBE4��c��=��3��bFڅ����,�g��v�2Y[[�"+��W�.w��_r�S��J	3��Y�H�?0V[9QkD�>�l�ܤ�_�����kp8CF-.��YW�����ux����"�T�Wr e�W*�}z4���3�=-�z���0���-�gj�&�aT*:���*^`�;�g��E~�E�1�J�:�$���s������"��A���p��KW�r�ХP�?�,_n0ps��'�F�-�1u�G{N�-U�d��}Y��2����"�춸.4�����,d�+
/��/2�H���-z#�����������4s����4��d�/.u< ՚�9�-ѫd�>��j%�Wv��Jr?]�8D��2��+
׺g7͂N����d�m`j���܄
������@�����á�1�d�`ɉ����Kk|����ϝ�ɀ� @9����9
����f����j��2���_�T��ԍoFΨ�^�<41��%[�M����e��8E�t~�p�H�Đ'1�2c����(���	^����ش
�(��Y'm����@�,�W����$�/6���:��KY�e{!��#f6N�sX���ު��us�4������/l��T���@w�1R�;Ȏ��CI����k�8*+zc�I���Ӵ�U�/��(�a�L�K��b�nii�x�L���q�I��f����_�:�j���W�}M��,�K�u���� 7<�~Kk����Y޽{WS�4K=��S�bvM�?���eS"��π[�	�Nr;��#z]�}y�k�u{����k�Y�,���VF|Q�&5wف*P*���0�Y�#�QGu(�(p,p��ͥ:�$��Q�u�C������sl)@w�T��S���U�1A\W:K+svυ����iW3TŽ? \�q�����g��L��ל;��j��E@�[f�Е�]s��
�@ƕW�W��E��{{{�Tz��ַ�����Ls( #Y>�P�\��Y.f��;xH\ZZI!_92�,�����j����Ο1%So���8̒� ]�I9h:K% �djo  y�*���qH�����̄�?�W��L�������S�M���E��x�����a�[<Xu������,����/�lF�䙡���F�pz��*޷�ٷdԸ�HL���k���� ����#}�)R����|���tu�wP��ѕ���⧾g�8�v
z�Ƞ�%H�ߤ4��Z880���{ׇ��[nVY�o ���J��8^�2�444�^�VX��޺k@ I��6U�� �_{���0)�n��
3x�R�,N�)�}F�Hr�TI���Dھ�W(]�b�XϚ�p��S�Ì|v�נ�Y��� #0�zH�T�H�P�eXɁ^P� 4
{�OPr��T��a�zc@�Vx��P�k���Y#��seďZp��w��#1ji{�S�=�AޓrAz���]�ior������`*�$��w��|Ũ�s*ڸ�~ꏗ��f`U�P���j2����g��kD��@*�8�Rș����H�Iw:YY]y�W�d隴EeAL����AH���.�{4���Y�o��RӞ���>Ɇ��5�{��$�X+e�ue�<Jo��w�w�UDop	����_��n�L��VN�p0�0x�`"/
o�7,ႩD��6�Z��$Mm�&*���:�����7�� G��n��t����l��pBҊ!�������0N�bڪ�1J�BI�o�l�R��{�gǾ��I?>��_��l�w��]]���f]]`G�N�n�}#�Z�8E�23�<�Ia9<�Eˇ�i��U���U"��ݎ�\Z�l� ���QB���z�������X ��
��`ޓ����S<Q11v�����99L!-�R���cb����z�^1���E�s��������=�U�l�\��ϟ�����(���t���r�y��3��~(�phg͜��A�O:�Q
9��]T%��
O���mr�Q�E}��E�m��":�4��B0U�:#@��_�Y�yOB�/��i�^
��� ���u��
�#n{�������/�P$�%QWW���,x������YρϚ��ο�#:[#�W~zpB�2{�C������go/|�6&��m�w/�X�Ei����b{4_�S׹�qlL����-5����cY \0�O_ }��zqQ�TT�w*.v ���.7�vhN������89�K%B��qr%��m?�����0C��8Ӹ�X���F��g=���������) �[���	�$2�j�&(���%!
�b��}	ޏ���~? S���0����B���'c��Ն���\�9��l�Ed�M��B��4��Q��V��9��B��.�Doy~�
8=�M��\ڳ��a��$D��x�W}�������45>'�#�kU���j�I��V J�"oQ7���𦚓ఔ���Q	&��dM�w��Ltʟ��4M�̌<����Lq$^6t�ތ66��3�c���j�
��u���¢w�&�բ��]�v��,@������Xh��-�]��O�c�K�(��&OB�ë ���@�E�j��R��כ�ƺyO��h"sx҆����^�\={Y�T-��5�T�$	�_��wY;�t��o>L�-�9�+O����.gȁ��v�=/*'�<��겊?:�z�uP�&��v�6�4mv�vb�t Pϖ���i�����ʥu͂��1��|�_��I�6ϊu�kjP�L1�����m--3}��	hJ��3�%�s �w�û��kLSAp=	aׂ(�&~��S@��=�����j&�2�.�4��P`00((E�U�Ȳ@KFv l~,�]��,u�n�IP���/̵�f�z6�� �:K+A��)���,���S�C}):g���;�{ar�ߌ�����wU�q���⠒ccjܡ�sB��
�cw2����a����m�d�g����wt�b���1O������y�=~�X���.�E�z:��0A�iW�t���X�UGA��Oxq�u����s�����5��#�@$991���.��R��&Vђ� ɡh�w�#�J	������X����(c����@#j�q���[�:�k5ת�W[k *�."���i���(�2Lb`��1v9�Q{D��=�J��W7}��h[����4���)Æ��Y�$%{@W	���/ kUV�����\;�8�sz�$H�S�M���)a�� n9ӳ�?c��,���a��4�ǭ�/ƤN}��)Y޺����'�f7X��r�ۣ��mIIg���]?�^����ҿ���dT�IY�M���Ʌ��n�C�ǲ����z�&\���C'�������	�"�Ȥl�ϟ�qq�!���甾/@�R�Q�mQ�eW��b��nTc뼆[��_��y�o�`�{-ӫ�s^/��)�X�A�æ��������r�έ˓�c��o�Js���HZV��]����P�X"��� �\q�U:A�3亂��8�����u`I�c�%�T��þU/ɚ]�F���1��ͻ�2��M�{�o�OFWi�N�M���c���rp0�8�@}g��� Â��UJ��R��^�����G�<J��Jɡ�K�rN��Vt�������]��[��JF;-��B�f�KK��UI'������^�Lgw������#:�-�A���4���p���E��#�=y�qs#�V�jƦw��{�p��Q �]��t󼜸uje���|qz���%i��NM�oh9]^+X�M�91��H�J�d4�n����Fδ�J��
5�j�d��K�?�	Ϸ�I{�w����8ch4��!N�F�f���m%#�&�h���%�.t0�.�_^fL�%G��/G{gBA�	�ĉ��G#PE�V���e�/55����F.іBỻ���$�|./i	�ј�;���˳EٵU`RD͓vR�q����	ҹ��('�"���;�	%P�|�g鉰��V��+���+���.� �+5Ռ3��7�{2������?}�/q&��]s�R�!��o�*è�@��@7���p����]�`.}�!�|m�M����7#D����B�C�4W�+ot��,VT	҃��K�����vκ}.qN��KJx1`7�,k�;�ag]1W�5@:~o���o�˝!�#�ց���@'m�:������%P���]c	�+Pk�T����MMh�j�d��;wLE蓭�+,R�/{��\�{i��{�6�{�%�"V782X@Ƶ?����Y��p�H�pNp�5�*���Һ�;�P�*V�9�=���'��z�+���\�{P���FQ��4�W���J��f�8�\���*[�jÍ���RiC�Ld�Y��1��ɔ�'A�h[�q��hԜ\v�؉�J���d|���vSQ����0x����l/I�J�'�� �7���BC˚1�X�=�Ajym-���F|��E�	(k�A�����F��zpdr���R�L�?������S0�q��(��͂t�R� 	�w��v��6*�ͬߦ��c'��RȎ:��˱;mh��
�*�DF��C�̓�^����"[5�+Lp۵t�=�����beu{�j����o�r)��@\�D����T��[�,��>	(~�{�2?2�$hR왨/]H�Iy��O�����V@
cؙ��������yD�G�,N��
�A�u��)@H�n�R�M�35���kE9_RI�R^n�b{kuL�'�h^+tu�+C�0貚�565̗���-R<@߃N~D���6v��Y��A}����u�N��hZ�L�3̋�( A�54�|��;���x����r~�QVY�]5���h-[��IǴ+�� ����'Ag�0Nbt$	(+h�f������-��:���?�	1?H���:��I�Fs%�։�޽�9���y�5�B�<�0���o�l�ۜY�c�1�_������C`�;	v_�d��	�b���:L����N<~fd���h^+��K>~~���1������d��}GU������<�
�0T�А�,���ɑO���a9����5�<�-��39F
i�?�Mf��C\J�D��'���/��7h�/���"NuǄ)��M�gĔ����}��	���MӮM��;��d��II"��K�P�4���'#~"�TJ��Cz�`���]�ڎt�q�tU�,b�>/�jÞ|O��&eD� A���J��c�J��9����1Hd�f�D�vG9�9��@B�F����ꢥ�g�m�/e�bT�ΌD4��|(;?/"}�7'�K�*�>'�O�
��ݭ
ޮY���U�5�]]_�G��u��
���:�hRV.�ǡ����O�I'�IF%�� KJV�*����I��=aq�� �JCC����
�>�vzۿ{�b�$.���ϯ��/x�@n�!z9��"'ϼ��:�|���)����բ_���)�a�aT���:gAm+ek��/��>j-��}�͆L�����Z�EP4h�I*�<3�t�2�7�)�K��?|����)���,4,5r�I�lÒ��.��J'�d��k�/d����A>�ABJ&�(��u���oJ4t>��r�S��-�ۺp`�

��l��Et�\�mcly��OO�+��--��?k`xηI/2>A�*s!�?W����,pd�w ��%��ea;����`��@�_	�����R�z��v0�'�2�g��7 �9@�����}��\t�aI����=4�w�L�Z�)tۭU=%lk$�:giR�r�t����Q��^���� ��~M�?N�J@TM�=P����N���)9�`�2�J�/�E��|_��*�HU��*ް�H����ߜu�=��W���}��K�AH�D�ɓ��O��{��"n�Ѕ6N/f�G��ԍ�\�_AۯC̬2@(��S+
������!㳲
 g�~��ʀ�;A����M���w<�֠y� ����$ؽ͙vJh�ʯ����zƑ���mYIO}��E߆��ҟ>⺊f6�=�B=w��O���Ks�7K�PՆ�'����\�j���lEt�Q\����eۚg���L��K���i-t�u89��o^'gKC���'��QhR��L]>�VI��Q#��s��*����Y���p���]ÊlYod���q2�oQ�=e8�ol�i�������]"kxt�fI7��nm��lF������D�ڴ�F���mKSi�}���rZ�,+�{�� 6���]jm]]���Z�{�Ғ�н���������E1���=����������̓���&����>�8nLQV5��4⿊�ȿ����ڻ��	_������'0��fQF�(l�e�=4`j;�|�2 _�L��\u��V��7�`��?ۙ_5,#���GK��i`>����nK�!S}�
���~��3f�Uuu
�-jjjb�g@Kr�L���N���?t�o��F$��A۞��u̹�����&��X�3�QMe�75=���3ڜ�E����=7�Y4��=<���Ws�򂐑��{��)"{����^:�ׁ���.�K"r��1��O�
�\�U���\F�S�eXU���Ǵ�����sRV����X�ձO�ֈ����I7ޔ+I����D�^��5ⷱ:l4,���q�b˯��-������ӛ��v��f=%ж�}˻�%�r�6�.�2_&�-�JZ4������Y(�%v�4� �5�)ʰs����* ���v d��!���H���_�u򵡎����芵��5�k@@��uk�I����@�O�����a����B/@�0��f�q.r?v���y�L��Ռw��L0��?{�����5DTV�r�'Zb`g����&�uW���Y҆��/����Ra�Ѷ��9tx�� Y�p0��hlP�}0,}�&���}:D��+`�̼H� p��l41𡃀  (�O��8�u�(Zߨ(*J*]>���u�؝k;��Z����jP'���u7��殪ި��>���Q�1���QA�9�ތd�Oہ��[�y�i8�%��g�ԯ�*�˟��*�b�~õ�~v���O��#a���%�~7��^Myt�)���	��h��Z��
�h��rt@�&��<iUO�����K���f�\A��us6���e�r�)����0hG�R��EY�}���
��)�[=n�9�Pr��ۮL=�-�QKS�P/U����������}|Y2�z�4��5�\����jG���S.��э� o�:��ù;}�ޝ �:<$�R���3fWɭ���~�tlmQ�m����{M�]{{$	|�w%���7< �~|��"����薋n��1�7����� EL�h��}utn.�@@:��O���G]]s	V���O�� ;��=w�6��XwO�X��@���3U�=�o0?&��A�r��x@�v[�o�p3�f��bgE&U��$(�TE�"@�E�Ղ�Ńm?~�Sc�x �5_-��HlN"�Ư���tLQB�R��)J2�gv��L���y~����nD��Z�����;q���Div�9Jd)I:ksf+p����131���	Sɳ��Ŭ�9����6��R�����)O2��B#~���{�݊G�k��Y�6��!M-�=�,��/*��n�7�Q��J�t6z⵭p���c�=��ҏι8Gռ�i8T?��J	�ȰVφTpM�>��!�
�<[L�!��>)|�t>�
	��fR�پU�ioU��@��ظ�:Z�b�@�ʦ�����B�,L�K@�RC��H_� F�F`߼�腓�oK�2f�yB�Ԏj��/�w�SJɿ ����9<WD�j��"�镕�|�7fa��^(k�V�/��$%z�|K�	 �DEEo���tY
:��%#�Y߳��"%g�k�s@��=��OO_��K��Hr�"p̀���L�]6)s�d7*���D.��n��&����DD�eZ@G��3V�mK��<˖���~�Y_��C<��P�˺2sXF�i`n_�n/�E��5�~���̤���zh�D�b��������#�2ktڭK�9�Op�+4��^�
���r�B���u����o�ju���a�Bi`e����C�����,�U�=pl��]��b����8�<:��.(%��kk���3ZP��d�Ak��
�Ά����X5KY�������S���;9�C���%^�+6�F��P[�̓�X��� ���j:�׻-�$* ���'�(��e��� r�����B���Լi����Tl��Z(�viD�Mz�\���,ʉP����vtX.�'����Ϡ�����4�r��н� ��w��xJ�E�?;_��č-@{�{���=]Yo�!"�Y�yw���}�o,���1��1��� m3Y�ux��}֡F��u��7q&�����1�FcU���y�kk_�ݾM�u�1q�87����«Ԋ�L,��O���x�2�E�O��PA��EYA��6�6!�r��2��|7��K8iѕdN ε~b�/0uW��ڦ/~ʣ�n����a�I��\�����8�L��f�^��Ȳ���tx��6���1����,��6$ض���D͝.fԀ'!W�/0�xS���bY�[<
$8�a�����سT����fM1�E�2l�������
;K0���B\#���B�`��끈|����
G�{��+B�����O.;��X޼�-sTV�u]�eyt��κRh�ӕ�') �P���r�"T����DD�]�}^�*��l3.�k��Aj�fxH���5�2��J�>�d��=�G�!r�g=̗��E^��~�	�Έ0O�0�ZU��]�M����؊¿���k��\��I.��8Ĥ,�W��pa��EOB!�&�������0kP5~Q�iJ���w� �7�C�����G� ?s���Ɵno��;&L��ǎPo�w 6ؠ���(��G�
;�˩DKh����3~5�zxx�zU��N�M�]~�%���~�*W[�m�JRx܎���F�u��)�k�h��@~�u�qp<f��z�[S�8:y��
 �D/����AZ�/ȺD�
�T+��0�T����9+�V���fP�N���!(�+N�޿��wA�+�b��%Y�Zot4������uN
bC�k9Д��v��[N�q������mTuAٔ�s�����tz#<F	����V�<ޡ�!5F�0���ɹ�vA��o�E/�̂�ɳȸGԢ���˳B�� ��~h)��#%�b������F2"Y�
�1�_��_��w����Sʱ�{�����U	C/�>��^Z��F��e�B�{n=��0h��=<9��ZŃ}KU��|Hr_���P�S�Ǳ� <4w���(��i�>�.��V���1H�4Tx�t`��VX@R�je�;H�t�F��J@���ɓ�Jd}�./�P�3�eRȃD�>ϧfݓ;^�g�8I/s�e#U|	���j��}cbbRi�a�<���)jA�#�OO��^k6��al��璒�}K��SU�V�b���g���7VF�Rari[�R�Ƿ7���lI�>�Ft��J�C��/&�G��׾�<d�;���vb��;����E#�9h[@��Xb�A��3�./I���� T#�����.��'M�@ٚ����#�Ts��ۦ���s�`�K���y>�$P���F�Ӛ�7\�:ʜ�@疞6iH�_�W{�)�L�e��^��j���X憢�s�"�V�X<d[���GlTSӞR���w�� .�%���e@�_k�J��\]���M��J�,��ʱo3�,���H)�?�[|�P��&&!����s5y@f�$�#��U��T�S�X�$�3�䣨���?�}  �EL�N��\�����������9�KA�ޭʲ��
�A��|K�<�v&�t�u rY�j�� Do]Y����ir��(|�_u�I}?�ѭ�CF>pN�]avě���	'.���7���/uJr���TY�L�xf	�db����z�2l�����O:���L�4*5P�Pkg��6oEE]�����X�2+B3+�Q?؜L쬷����S�$44��p �O��	^�@#���ϼs8 Z����&�ս�||J�S[{�[m=�$W�]���5�㣩����@���H���1nZ��H��HyP:��E����jH�	��1'a�c2�K������ t�k�P�\U��U��6�:��#����z�^v�3#fSD2P��7�.�P�?��� ��S;�?C�C��KM}̓B�5:��I�/�|h�jWϝq ��S���@I�{qs�߻��j�����cwL���/��܊Z�����ɧ|4@�^m���>�v�!{���m9���w��w�USJH X�|�A Kޓ��56Q=�H�$��ԙ �0�.�<���]��@L�m䵋�� ��U�3��@mZ�UA���{���eM:��w��XK�Nb_-A�F�X[ձ�����aB�G\�#MC�_�іע����t��<b��|*�;!|�|	��!�\����|��؀VI�)"=<�JCN���P>36�������VB0T��ms�fy�ƹ���9{�Za��8S��V�\�W�zh�Oc���ny�	�ɺkqx�	9���
�sv�H[袡���c�	g�2Sd��&e;%zx��ز�^��t?@��S揫8�k��
h{�ڔ� �$t�0��S�1���.��w �@�
�RO�
�c��4BfP Z!+*26�u�P�[� �����S��¡�m�S8�Y����ָ^,�D���ja�sIŦ�u�_�|�hУ|xCgu+�a�Ȥ!(�I�6���� �kcM��q�S��.�_��r�	���+2q�����9�5n��M���|�����.t��4�oW�J���:��N�9֋wQ���=FY9����5�AAqzŗ�E���u�0��,���sYl1x���P�����I֗�v<4���owU@W��B�Y��պ��w��������Rx���.���7�t����7�:~,��p˭~���!~'[�rĺ��6u�� ���%;A���1��~e���뒜j�'[�<�z$���ɩuk~X7�k�$KGggi���{��9=R��4蘟w^���E��<)N�.�ɯ���LΆ'i w3X�Ʃ�����[xx\�:���/�C�PON�S�\R���y=d/���h 5�U����z�(���R�.�����
HHJ9��t�HI����R" "�0CJ)�w�������r�Yf��>�{?�w��
vk8TV�ʩ���t��ftx�����,�[
N�� } #��$|g�Ĭ���r�c)ly��2�أ��6=��pΔL��m�$�GS�ߋU)��i�)��T$r��[�_$c���eΐ�.��i|����[]��1��.R@g���
BɃK�j��������H�>A�;ff7F�N6�y-�7��X������4��3e���<A�l��Ѯ�� �j��f���o�G�0�_�vLW������Q�V@aK�k�T�|�ᶛ)�@.X&���N���ѡݹ� �6�v!�!�I���-�s��ܩ���k���/j����+5�k��n��Zq����;���ds3G�׽9����+���i��2��o�?
����G}گ��se��= M�o�Z��f?n�����r�o�X��;���{�����H;QX��Ύd[��}���d��pm4�3�����1�J���wʔAZ�;����n>߅<g�S��9z���W��](������8���/-����
G0�8�D�.gqH��m��U�ɰJ�P_�5j�w	�||�T����c"@h��'=!�5%ހm���7�\��b~�����X���a�V���2�QD��JǇ&د%�D�t�A��۫��fF�MY�=�j@}�e�NN��*6nF�8��1S�Ő�d�G�#��ˀ�*�T^/��F�d��<�����8 ��q��Z2���+O呕4\�����O�&������ɶ��:��� ������8:2�-�߬����<�r��9!-@J�mRq�\~B��z
S[��Ӻut�{z��V��:��ٯʘ�;٘ݘ��]{�l��d�����}R��7���B�$���R	)k C�2��8��X$��]�!�C_}��?�'6N7�*[����m�e�P���Y��՟]�����k�g�r�(�j�r��_%.��M
·�Z|��$^0ίR���Q��w�ٽc�R�ó s�����&� �͖��v�[jJ���Y��Z�����)-��T@iV�ܣ��~~Y����>r\j���s��̪�c2�e�c��2�p�n/�O�ڗ�U��M�'�Ky�*==]Q�>�	<ds���n׵��*~T	��ME�$�<j�h)-M�����2������EX��C`�S�o�$� �Fv[&<QT���"��K�<ї�	r��`��\$��f�#D��ߥ���HAV?���\�5k�5V�p�:����E���9I����v�
;���3�������p ���j�����VVV>��L(J�juO�)x-��0�^�KaqH�t$+�9n���r�=Eo�Em%F䌅"��ᴷ�UA�&��tq��#]�z�!ul��U�b1 ߿-퀘~�UBSV�)vl��Y^N�c�JI��߄e��˻�{o56������}Ƥ�[l)����rd���q�d��9q���_x��eh0������D[�1�<�]kt�ѿ��/��l����M}о0C�.���F����
ʣn��W�E���9�[#S�R����َC-i��*����&��O���%V��#JK�����ȫ�4��_���_��Ѝؾ�s����:n�~����l�J_�+Ji#��8Q�;k"&���Xx�^w|�� �o��Q��BP�Hr�c�"n~���AWW�&
��	B{8jobq�/w`}0�����dO��T·�����<<�Nl�U���5ߪ�:�;̴�M�����3��]����:��@Zh��Q9�4��d��*-��q�lj��_f��,���Ϭ����4��ci�=Gk"�u��퍾�Lo�������⌎x���3��_�>��Π� )��u������ҏ˲���� ns�ׄ��t1����-��!q��=��BQ��GGJ@d"3����C!de媡��1����~w�?�h&�&E,��G����m����M@��fM s��Ng�s�:%������ڭ�o<��ee��ml �%�� z~�6�p8"V���h@���[瞯���滈�_��r��� �pk,'�S#����\��!��k@��� xc��L��-���6P���RiiҾРl<����B��4�<匋D:�.���wp�0;��l��f��Ⱥ����EtY/��@�М��h���Ғ��������w����o�w�_A:8ˁ
�F�ffpp�����&|��ƍ�:����r�Y@'�k~�_�[�A�VIhE�];
.����us9]�~c o��q�>�)�D�
����y�)�NMz~��\d�͂o��hph*ڣZ� ���	����z�)<�eS�>=���6L\���C�@���B�I��|\j�u>ݾ�Wh��Ӛ�𒎈 Q�$�M/1� ��B2��Ǒ5���Np�|�XX=�V�k��v򆍈�������J8����щ��=qs2w�p����V1�0�]hx�[�(K�Y��ۨ�ZZx�I���P���{�k�Ѧ�R�ԥ�_o����͚��u�%5��]�h${[
3��/��J䲧&�����bh���@���S�3�:ԉT&��FfOD��C~9J�P�~��^|�D��'k�qqZ�ͫ��̓�1'7�e|hp2�&�4���(��v�m�X;���*�pKKٲZ��o�cPű�����\;��Ԋ��>(��݋�����˥�?�5E�/�+-=\-���=r7��8���I�S�d�}n�>�Wv�����1G������:�c������W���>hj�e0!�}6��8ܾWT���w8F`W(&&�4���B^'�����V�����Mfbjj��9゛��@��$��p�c���M
�QǪ�ue�D9Ą|E~ɠ�G��rn/}��g'D�u��X� �L�w����mo���|�y����.�n'J��r����*m���p.7���FȸJp�O���������C�R�um�u-?������~�#�9��{⵩�~���)"[���"B<ى癿?��zn�)Cc�X㷶 }��k��GT�����s�{����ZU���QG�����\T���W���������Yn�y�U;ق<�7[��fB�AOZf �!-���a��_+���m��X�ҫ��9���<1!�C�
¢��@ s+��su��=��'�z�^�C��Y�CW��	���o}�����ӌ���m4T��Ws*.�y�=�p62}X��<�F|�S������hDt�2�!{|m���}����4�b��|}�[n?��)��%������#�h�<��KҀ��ʨ�'O�eɱ��i�G�fEB�z�����:�"��3j�<Wu>[���)��u�G���{���z|�Jx@�}V�_���U@%�ra�k	/1���̠I��G=��8�ԅ6���w(L���`�bY�x��C��#Wl�=֊��]�A(��k�(�L�RM5��u*�_7���Aw�<��	_{��<�}~������c1��,Yv��l��4t�{���"�j��}��nB��@��2)�JE.��n|��Q�l=�4'Ue�pޘ��ࢢ[H��y�ҪkkÝ`$A����m�W�ۻ�'fm2(�͙��P��x��������OS�%��������0.�9�y��2��t�{�q.ք�q���A%[�ڎW� C�$Xp$b��,j*�{랄Ն?ܬx�I6WMF�i��LQ^�śڗ�V�g���߸���*�:�(EȌ��fE�أ�{�3������4���O=�GK�}��X�����q�8௴������^6�Y_�V�	�u �R�2.i@h5
3����7oȇ�=#o@�z7��@����:ܺ~4bk��5�T~�1��)'��|	&^�XWa^�!?u�1�;��|A ����FB&օΘb8���\t�׀E��N��nP��`�rr�$��*��� �8t�z���|���_��ڛ��_�d�=8c�A��~T(��?��wI)
��d���啕�'�k"�����k�qs��ww_IӚ��·oV?�J��_113����Ԓ>5]i1����v
���q��wu��]��w$B�p)��2`K��	�R	7�=p�cy$~�zl5��)��#^��S����j� �L�M�fb�$L��.�	4�|�;���.�XƜ%�p����Aو�L����Z���a�|��B,)�E��]�����q70������\1s�C�Û�z|ፍWpJn�;�X��������.r[=���S��W���kۼ�8g�w�`�jRX�=��/���#*w>�*p�p�`f_6��v�������.]?^B����բzI2�u��ݽK�DME5,��� / م�]�����r�;�e��L\�u�O(��@>��ө0 TV���1E~u�������dlL�Y�GX��-�\6%]`�q��$s`��L�C�B�B���k����a�����)����]�*�7��v���%� ��ϥ3[x��7e4�7���0�l�o�O�Ă9썑N0h�g�+��--x�ӧbhAҵ5����^��������g����,��ݯT
$'����%500��ev����.+�Z��s�A��N��������C�]?:�d4�p�ꜯ��QDv���Ӏ�T��}�C���#�6�(�^b�����o���vf������/��w�s�zIY(�>sG�;�e�q��q��0��׸,i�,��Xd?��'�v�*^�[I~�1l��a�[�j\ɋ����n|���Q����3�H�K�3U�[HL��5����� T�7l����F�]ֿ�{_G���#�*WR�t�` 6�`��H*"�.�<e�B�Y_�
�}
_�����Q�W���k�-E��W0L�w�@�ݱ��@�pP�k����eQ.7(�o��I�f� 1�ߙ�hVE���B�K{�zx����*yј&C�D�m9\����]�iG`��/�N�e^����S��o�oK���m� �+��4��/=��vln��O��^�z��ys��՟?[��d��=<�V�����!�!.<���|j�@>�zC����4���� ެ�N*��	IP���vc��8���cm�,|�\�R�/%2;�%�D��
E��xa�C�gYM�}Ax|�<����y�5��6�%�>3Hew‸�@���&��)	���A�;Hw�1{X��0�36q%�.�_MB�Ç��@'+~��8- �&@�>�v�UFD��I��6J�%��U5 �J�6�/_�
k &H�-����>����d�O���c�����1���. �CHx_�#��>F��11���ޤT���!145�&ڷ"�����Ąb��bw\�n�����ov0��׷���K�o�[(^��9b`jJ�8<Ħ�7��|:�w�����A��T744L:"��m��&@l6|��ر>�q�Y�H돫���f�JN���F�=��,��G4����x�m��eX�{�qY@|3��o{!_;�g��ϟ[�H��a��� K�ګ%�����rFĲE���}��\,%--_m��2'b�;�~y��'"�'�Nk��^m���22�[����\���(�3o�?�!�ӧO?�I� ��GL4��E@���j��[c�*א��L�|.k� �h��ꬻ����.��O�?�B��,�!�@�NOZ������� �Љ��dk�r8(J����Z���)�rx~{nu�W���B3ZY�!���e?������m ����(;��_��ۼ$����[��������;��8ɫ��"22o�'����G�e��'''�"'0{�<!��_�|IZ����y	S�u��f�����}���.��K]J�)���Jה��J����U1G�٣`�C|"�P�v�<!��o6��{�=�֨�O7fr��5.Q����]ܼ�LN�f��M���r7}e�����Z2&!�^oMY,��A�������6R�[i��B9զ���o��v�i.�ŞtܾlG�*B�2�f���l�?��W#�%�Qj�oi;i�`WU���Y�W�~dk����o̞K�Oe�}5�G-8�����o���̪��U#��W�"���-���"���f��ζ��}(��'(��L2x��8����@��CE�]ŷ�6~;(Ւ*Y���6A�����
���X��e'Zγ_V7L�_B��fW��o*�	�I��u%ف��ٶ��bBB�����1�~)$R$o�fV����%�Y�k���3Su�=��%��T\�rL�����M��.r�R/�'�./_b�@���ӏ�ŵ5���h":::�\9@����%���e�3�-|OĚL+�?�tR����bFōD2�k��J�Ԥ &���_iz�D� �"�<����{{��������b��{���F�&��0����VX�A�XV���8|�4�>�� �rҮON>;G~v�v��P�$Ƴ��8��d�(G_?q����~�J�Z%�n����:̡�4�/*WFӹ�����4��-K�}�?�R�w��V�`{���Tb�׶3ƌ��|",fvw�!�e��
�뻍�4���v�z�j1 �[dr2��$�7OY�q���������ڂ�&^626�y&��1�^����H��1�j��>cv^^p ,*|ိ[���Zi+i����'�[(���m��P���}u���⥦=�qq!y<GT����U9av� �DE����=����^+��2S����&6��^���k��?�����C=�Zޡ%Ξ��Ŧ�h:K�p�Q ���O�ޘoQ��41�O���N����1��
@B�8�=��U�굯���3�yP{��Fөb7T��фne��,zy	[�x_�V����,���Cž�����ag��4��
���E������\}����f����AlQ�S@��B�����=��%`@I�3GC+�Dɚ* T5��a��4�D�� H�%E�V�����%eX'�.؍~2�PiC��՝�zU������'�y������8���b�ru�`z�~N��uP��u���Ο��7U���PV���H�5 n������k��JF�4��iI�z����Du�-�������{�ӽ��kNU����g�Ƭ95��c�ۊxO�Ͻ��ُ4ܧ�%�L��˔�'#@1r~MzXc��h/����&��ft��l0�/2��ur{���66�P�I�h�q!����������w4I�LE�rrb�K+���C��/{^�l��ܳ���7x�+;/�`�~1��9G��;��L��p0������]///���F�+G0�92��n�L��C�'j�K���r��l��rx,ɠ�ig'.���V���ur+��f-����� �߱��^RAe�}��D�E�2mg�?FBt�İ?`��G�f��Ȝ�+��	ܻ�AQz3b��tb�Zة�-�)�����^a@��I����D�`�c�$f��#�.��\w�z{[�',n������ň���L�倿��'k@�F�epF��L��?|l�����J�D/A�X
,�S|(%.A^I�
Ǘ=YX���I
�E�@2��牯�]@luƚ`}�&^��q����-R@m����DDuw�"�Å�*؀�VTV>m�����5�1H�g|ʑ(Z����Tm(W1��O��@���7�t�\[#�2\*j�|�X�T�� 6�%c2�4�=�d�Iخ )��q&�@ 9Ȃ�%����/p|_�8����k;�v���4Z����j8���}��晙���j�[p�#��[���F������A]-���ל� L�ܦP��f�1��j���8ς^�o���T0f=�*�'��wTo���G�(.C6o��m���a|W4�	ɀm���"�/Q2�J��041	�"�\�΢ݱ�c��L�����v�фHe���s���J���r��T��A+�v�٥1�mG��*��P�C��nE����gS�MLL��+]x�����:coR�7�p�����BJ��r�Iti�yX��(�z�֦�4_w#�7�B��6o���'V�����/��q5i��$G)�����8X�X��"��]�o��E��R�+��苡�1gg�Y��� .��B��������W�yP��N���ǜ,1bp�����n��+$Ȅ�j��^�b_��A�Ȩ�K1�
�,W���]���_�?��ȥ���TxiCP�3	5s���jo�N4a`����tR�j������n�o��r�ջG�����WX����ZoD��� G?1�<`�:!fs`˅��}46�t�wt�	�2�����U�J0-{6���9��f�(3��k<����,O�������#���ͱ�5�N�=y�˾b{�w�9�͎�ȝ�=U�C�հ#]$�����Lv����C����1��!.�gT�*�9��t���cJ2�o:(1'ggׁS��o� "zX�e"���w;��&�JJ���Xz��EDj�W���N4Fn�s�#m��P�c�W�4P�Q�V�ܽBbbq�۴_f��W�ڄ���I#M���;C/y�]��3?��8y}}Z���{���l��8�b6�UR,��f��s�s�/7Y��a�$z�����<%%�s1n��_1�l�!��iii3��'H8�*6n���@��a��G8�_�� |�q�lj�+1�����eUlDg%�C<��Z:U���\)e�fgg�{4���|�'��Ϗ�8�8����9�
=����� ��.��c�,\���;O���9|{	�ڃ�~���� g��}Wƨ�� Ui����ss;''��^��|F���P(�+K��@I@;����m�)x俓3��}#Rk*�FՆ��f
LB9ܧ�ু�;�!nf1�}���:�_�;��G�3��uQMNZN���#���"iʭ���B2�	q�8\����+X;��\�H��[�'.�a]gQ�Iaeݸ��@��g5|��1@3���6��c�	��oqc��W���Z0�?H����^���gFL_l Z�U��	�?e�L����t��{��FB ��d?*�\�+�g&M����}����Ȩ�Q~�2I������������9���O��=I&&&�7Tc؈���P0���]y_�~q��t�c 3>-�L;��~�:\/q(DÁ�}�\���+�'Xn"����ݕҥ�/]� W���b�����{�z��*O+r�/:6)H'M��KB��h�\�u{H[M&OA���t�^�0^0��\���qo�ZEpݗ(�Q0R��緕�ݵ�3{|��XO�lDHF.ԍ-+���1��tx�;m�e�D����̽lg��<��B�C�周f���������罰�/Xۤ.���%�' ����;���8�3�Z��2̺eh:4�<���~���	� �`�Ŭ�/ވ��32RO�,"�S{{�Y<2r�>��Z�v ��Y�`���|R��h���~��KM����b�^���y���[�Iн�*��#��Ԛ�܈�+�/@����|����K+%��$tigN�/�sM�N���Ƿ�i�����l��PRr�9�=��)��˾z��eO̡t��ݽ�$Sw�ލ�Y�15�	u�� �77?pr��>�&���W��)_�C��y[U����@	%��h��+y�t͙���5#c�Ml�a�ׄ?�7tMB���E�L�+
�a�ڏs�}7qS���.//�c
N�ʔl������'n���z}�ݠx�%Wd:' ~ȶ��N��ɗ���	Ω?,����&�eБ5,lJ���ۿ��s������T����Ib�u����>��T+~�t��n�Ie��xK,�]y|�OSp��Hb-�M��,����!�͚g�9.T�Ƌ �D��*�J���-f=W�ua�'�oq�ѩ�H���"�+m����*�.�� ��{ו���N�$$%�>��)�X�|����o�ha�_�+�ƽŭ��j`Z��H$*NWK	**��;�c}gOq������/��l%�� ����V��NS3�g���v�\||2�6�a�C�E�~>��d�lAOn�z1G�,]Z������3_�xm�A����Gf�3�K�6�2�f�?D��tRWrIG'�x̉��Q�B��e��?8��0� �a���F�g<�R<[�� ������W��@��HQ�����HI!#J��7�Y���f�2�[�b����AE|��$����JET�ah�W	�ZZ��K���B�Q)�w>�w�p�z^�[c�e54Š���k�δ��*�U�Y�׻M���P�®:m�_���`�ퟲ?H
	E����FR�����Za��x?��)��nT�b�sW_zf�";u֮�������C�s\����t{��(����'AR,�h���_��\�&(\�'��6�X�pÍXF�\�ѣB�W���9:��J=)h�� A:�Y7#�<�4S<�C��q�	��~�ɴۘ���]K�țGT�����
{�� df�~k<�4��uӰz
��^�`���̳���YcG'^�*��N�OK��V��W�;�=�ܺ�=��]��F�����~�AY8v�L�eu�V�t��b�X?������T��j"�텴��$�#� V�KG��W�nk��Od�;`��m9\�n]4�>��E��)���+��Ȅ�E_>��֦���`�R+�ҥ��K���55H���Ygkhj�v�,��`���~��w(�2ɫ�E_���v���G�]�s D�&ܶ�o;���:�N�L4�������������W��$$$[G~��5P�l�鵋/5��21X��(x�E�R=.� �{y�lR<{��F��qf����K��������Y9	���_���pN��61���d}QN�%8���KI\�XU��P�_�������&y6K��z�M�)s*0�x��3Ym��7n|n,��N��;J�$����$.�V [:�����7H�}�U���m��U�"!<4��K-��Ʈ��@{���|��d�⏒R� l�r�Y|�K�r�+~t�o���@��;{@ɼ�O9�����e��Pҝ98`U|W��}Ax��
]�<��z`���Jcm$��t~Y�+-��"�P������������MQ���{,�y��G�����zO�Y�� ;��2 �X���%٘J��Q���`C'�__�uX��++W��wh��W=L{��q��&$S���<���V��I���oQ����C1�W���!��B�8&�7Z�X�dX�Ym1�gm��nք�� ?�+PR�x�:|��3YR�?v��C�]cF��`���-
/)OꉋdNz͟��jԣ(�u��;f��r �9@����ń��_iyU��J�饫k������!9@@,���X���n������vihk�͍�<����ʥ��u:�W �B���A�v�| p�±��E3����������7�U" �}a�� ѫ�����䃓�����+������a��0�%{=%ʛ7��`�/�5T����j���������8v�ŀ���"�M�"��KZ�<��g����Â�>��B�v��	}~�l�\kYѶ�B��}n����?���=޲:�a>��R0�ϟ���Um=��M+��Y�����2�eq���ەy�����ʼ=��Pah��¶��V����}�k��]C�n��8����s{�푝Q8"Q�y�ƾ�g��
['������e�����:���6���mV�苛A$r��:������%��~UD�VL����7��2�˃���|�(~�宀@��a�r�N������Ώ��j�G5����SFG�����|�C��䡀��d����R^Yi���7�y;E�ϸO�m�A��l��V��ss��cRV.�Ý�@���v�����dg�t��\O6!@�A�@M�1�0��_4�b�I���w;�Đ~?��|����)=c���5�^ˇ	�d�����de��釣0�˾R, c�å��q���|��er%�� ��[���5��@9�h���0�E,���B��D`ܾm؎��3J��/���(��ؠL�.v�<�V[~�$���l7�ᗗ7��T��¤���»��λ>��6NK�!!=K�Up2�s�=�J�C2缓@��2%E�C���K���tY��=��ϊl�gGFn	ܻ礮J�Dh�66���\��o|,�L`|Ni���M�3;�--��,����n�� e�d*��,7��Ȟ���w޿� ��4u�����\����x�5��#T !+� �U/
�#H"�����"��S����_.�D^=}%�����i�K����o1���n�,�͗��D 9�ܻ�q�l�:q�OF֧��t$Fs��G��R,�of\$��Sū����c��vKq�i*tb=�y�,
|�L��qXz�EwOD������ݖ�����14M��zv�'	��*G�/�k3�/��˓_�lV�hV��द��n|�ՃV����`��=�BB�Əy�n���Btw��9�E�l�������;����ik��?j$����iȒ�Y;�4��2M�}89qvqu��k���;�mii�GB����$�ܿ�0��[��0`���������]3�_:B̨j�܄X�c�w$UY)��e^h\Q��W�U�V#�^���1|b���B�1����z��8��A��L䘧>�a��qWy(dݚ*�6-,چ�f��/FJ'Uw��#�W�Q�0^��ѭ08l�f7+fW�r����9�g���V)�90�]���g�߈Y�&B�v�{�=�_�=���@iARN��v��d�C�/%�3��!�3�3���3��ȯu��=ր�b��9O_AYY�ڬ+ckd�UU�${���d��NW�x{��|F��CB�*V8~�mI�g���ҠJ���ߊ�c�uDȢۨ�x���?��G	�B���ܟ>}
[Y�I�'�o_Ѯ�=,��ԜxƇ�A`��*�Y�oVU��;s|L|��oJ�&�J�n���[�� %{z�r%�_��4#�����H#��>%��!����"6(��N�~�g#�R����sں'Wg|�7/�j3�	��"��Ӝ�6'�i~�k����Q5�h<��Ƶ���(_�;�R�S�=��n�7-��C�&%�"(G��z:/���`6�!bsp����vCN"K�WIIv��{���T+^P�-��z_��%�ͬ��I\�!wrr2�ћ�����������;�Vܷ�����4��,\]�gV�Rԯ<}:��CM���=�xv%�sV�~Z�����&!��R�Y�D!�g�!ߐ��'i��-^lD_t�n�% Ǘr,1֊��}�Z���29xb]����"�}�h�'���0���^�DR�g���.�$`�|�5
�/C��ҹ\jP�#-1��sƓ������	�C	.�̞��0{X=+��I�w�@V��T�Kr(�ݒV��[u%dEo��j���<*ݡVxT�r�+�\�f�yՀC�^YՌ��z����uq��lZV�� ?�8���}3�?�GnLP�Lk��$b�{ٿ\Z��"U�,�	~��T3��02>�dS[[��X[������
X^�@m �h�s��D]�+���ѥn�u3A�
3_�i*��ttwEF�{�X�=��[��������=@��҇�ݾghMO�"nʸ��C������Wk��B��	Jx���������ʗB�u�K4akDXV�k;o�-���r�@��� ��_V�p�C}���+�4
��hۧx
肍2�a����wb�������o5N�)��{P�s}[<c�խ�81i`�Y.�i��>Vb�W�.���ey.��c��l;ٯ�f�{o[�t�4ɔNm���k������Q �3W�b���+���0UY������'��rSӁ���4�Xʚ���R����FFJ%<�L�D�/�d`�g]b
&O�KF8�>A7� �4��j\��������A����i�XV����ˬ 7q8;^��U��<�]�#Q���]�@I�*��_n�K5@!96����y�	&�Wl�t�Z<-f�]׾�r;U��:.����t��J�*�m��w�uω]�(6"J��QjU%�qo${
�Ԅ�ˍ���?z�J�-X�<8Рk$-t&\��on;B��.k�(����bV6�B���}ڬ�:WW3W�>�UE�;{6Oڂ���/�Q��N���n����;z��k>�0<<�:�h%պ;����pGFCI.("��}���IIX�9���}q.M��<�Ŋ�#b��.����?����J��ޤ[�*Z1Q]�c�M)Zg,ū���J2J���i��G;��mJ"i�#?�j��t��Y���9������)��s\/�n}=�8��ס*'��u�0F�z������0t�ڶ���G�c��ԗ��4�My��Z0a��$�b�xl��ݿ�a�sz-��K3pS�q��0�y���VwOr�c@��b ޠڎ[>S��C�ʎS����nS�323?KE��{V��0�S|:�`8�Խ��OmGo"p&��;�C����16y�L����&�A�'�[�r�I_��l`����5;�+�!
C�6�^�=���--rᕌ.��Qsg� �̪nD+��YS'q�8T�q��q8�89���.���|�n�Rm('���/��\E��hM'u���7���Pj� %[��6e� iWP%��)�� ��ZE��V�5�?,7��U/r��+(�/�+V�ӽ��`a%�$�i��A�\�S��m/��^;h�.(�ԁ����`A���++N���j���΂[�:k�v4�*�������7+�����N�ґR��R�kk$�M �rr^��H?&*{Eܙ�hP�}v�@4+���pI��૥Џ�� �g�x���G�$����rk�,0�ʟ�Kp�Nj|ߣ��yݷ�')\׀�/�<AR�[�@3{o (�PK�M+o�:�P��@Tl<EL(UtA�������ط岏>;r�@��p[����O+�a�M̝��:�v���2�A���EL��b����t�$�k�&?�l�a���Ɂ����g�'�ퟞݿ�
_oS�q�I���V�K6�J�������ihb�9[�t]R���?��3m��'��ܦ��� 	�H(�ʬ�<����N4bo�L�)T�����s!j��KZ�Ǐ�����U�,�uZ'���#& �r�~������A ����zx�3����jb� 0�WK+�g��I$�E��[׊c�@Nלﻌ�c��k�����h o._�g�e7��Ł[Yp����ae����C A��MhI��C�.|"�!���y\j�e?�N�qt�e^m��0�<E�;��������v���.��!�.z9���^��UnS2��U++ī��̀~n�ߚ���؎1�vVK�K;VSu��v3��Ŋ������SF����
)��Z\]j�]S���olr�G=���~ʰsM�i/���P��%z�Κ�L��[R��sD� �ӵ���'&��3y6�߻�V���Z��ߜUmH��MM3o�֑=�6;-�<�C�Aӥ��B~B�=Q�C��Pyդ0�j��֢�#W :A7R?��i����$]Y��Qv�h��Ika{3�OF��rL��'������k2&Kk�)�C�|�޿�32R�1*W@׽c!ë&W��6��W���Û�V���.��B���N�t���c� ���ǂ�穚͛S9�f�\���w���.��|�?�=����<���qu�<姶sj�*T���2Α�T���4�v!./_b�xA�����{KIX��h��D�Y���J	�H��o��b�],Ñ444� *�wi�>pK�^q�cT�O��v�X��A��@��N�hc�}<�vY���ݘx= ��Y��{ ����.���]a��F)���1	�0N�S� D��@�➗v㤡��B�׋�q��Ƶ���x�7m�Y�E�%���&�&���4A����k\ޤ��ש�m�p��Z�u�Zq��oR?�cOp0���>����`zӆ�����/nU�B3A~r�5�i�a㮸V߾�>�Sɝ$s�g��4!}�)��fT1���~�5��; J����Y�M�@l�v���7UG��+a���c�7-���===��9��K;~~�u:��s壗�22��Q� ��_��5�+.�堦�''h~���������f�2L���r ���d�'����>�9���Y<{z�DHx�g|��ѫ7J�z��GG6վ�.�39	�_�`V..�]]][�-v���?
��W���m:>����X��e�N��{0/--E)[�
���l4��0���[���+J:*�����%��@Z�<C3j��H{��=u@�Q��U��+�ŝ��Q/,�<z��m8f-5�����6�RX���=%���o�A��R�n�{{���Đ����6���k��{��~�3I$"��כ*Ƒ�MĐ��#�g��F����A��u�razz���;t����V�Zy�� ���\M�U�|O�$�`x���}a��o22n����Z��~H(�|��&�g/_��^�M�:�h5S�e)�(V�v[6n�*����H��<T������Y&��5��31���k��;S/��Öxl�5p�_ǌ27���(n��J�9S�������%��^�ȽzuR��Ow+��4t�6�Yo�Yqg���"��C{Efzƴw�d��qCU!Ƈ�#���O����D�e�idf�cN%)�Lw�e�է@K��x��O�����<�a�����^�GtmR�>�z^{���4Q8&23憆a#�+H�� �{=������5�7k�[&�<ʳ���pw�M���Qp�v_�l�b�β��i�����Ѓ�\xY���@A�W
^h"��2z��{PTS��DY�?���vݓѳY���Q�m-XV�D�'4�_���������Gf��Hߕm�Ev˱m=N|pq����J���9 ��~������T]9*9����`!s�6]����{��+�]�ٻ�k�t*��Fp�s+(t�jd�h�A�Վ)J05�+�S�9}A]�պv쳾�)�NV�ƃ���3��GȺ7)P�[/��w���q4]�lf� ���K�D�Lc�{��O��UçOm�qqq���$(@8NN�o����}q�~ci�)"%e�����<C~:~�f� ��z[+H��L$����B2���/�N���?���3Ԍ�zzAW��q�,"?��:r¯NO�"�q�v�r�Ɯzff�""#gݛt�F����J�~���Ҍ6�L�[#��Q���.�6	==}GGG�Kr%��K+ ��[u����f�rz�Ҕj��ݔ���M�]Y�����|�yV�XI�B���n��u��u�ؔ��
�>�?���v5Rt=PHJ.��]�,L�9��_��\�+]W�&�O�{�]�����32��I��4Y��/����Ĩ윜���N�^m�/q1ۻ����ѧ�Jf���xSt���y����ۮ��{M>��3ss@��9l?x]9��͍X;O&�iv���v��h:�x*����B��!���#�Yɱ���cdfo�압d{&!�ӡc�8f��]����?y��u�������k���m�Jԧ)����"��yw�<�{�8��k����w�ֲFuR���DH�1T��������R�lT���N����C��f��X�ʾ�j5�,k���2�@�H�M�W�ډ�-d�z��Ӣ�y�g�|��]8��Iĵ;��P�Sa��sqi�Jk�a��]�W��u��JZҋt�9՜�����@VX�$�"�e��E""�&m����h�[�##���34�Ty��	4�y`}M4\H�uE����n��!D�m߾񇇇�㆗�nl0��i6؏P~Q�fl��I�+��,�ֶ�ʦ��#**�{,�=�Z'��ח���W����o������IIt��鮸ջ��θq�Dqё�M�s�����*߻)3Ʊ峩p+~:��	u�����i����ӫB�Sc^�.v�o��B�����t�N%�RYt���+�q��V%=ŠKoP�θ!��<)9S4�=�����	f��.Q�7����;Da\k��<F��9m���k[;�Sn�pYG`p��Ke��,%V�d9�R��z�<����afe�z9=�t$����:�LŮ��(�(b��Q�BaΠh~�26-��n� D3F�oA��hu��F�-���G���?UTl)>��2�@���6p9�Q#f��]�f���_����J\Gj�A������:��ƥ���
��n���xE��Ot����I��h��Z��@����ß
m����*3�'���K��p&u�yh��Y�vfvvB}���%3��8���f�̄X8�>?�^��e/�B�h	T�"�V�p�����dy�������ȗ�Vh�%�m�8��4�2�}�[ƽ��o_U��<��0�Հ�
����+(�a�O#��a�H@O�үyN�&d��u���l>�\'�@��\S5Ӵ�X�fSh�0�sM���2��ۣȾ��������O��^B��㝔i`�������@����Дd�ۢHeKK���M:��_:p����B�f�i�^�����]^P��/)2_:Z8e�7X�GEF�y�p�]$E��R���b1E˔�����宮0ꪢ����Ծ��q�v�]6�©�E�S����_嫪���nlZ�Ԗ��p%Fn~ 0s-�N�?'�ᄜ�Ǵ�!�D��jо�����.|�Lj|mo
���TM�6��k��`l�K�T�M<����̫[Zz��	�#��Xht7��e����.������h���+�&<�ƻ,��0�QvAA��w������v�a=�e��C"��W3M���H��j�{�,[[���"c��wɑ��& �!��Sh��$-7n����ù�1���?B�Fk�C���AoRp����^9�dB3�MOrt��̘��������}�|�٭�͍����Y�/|^�u�.��m�>ZT����QP(���uJ�2�K�HRSD��H�s8���q�@=[��v����!��!��v�*����!�%������V���*�luo �-��*�{�b��GoC���keP�	*	�!~l�1��������k�T��_ut�薹)f�,5L{{yED5��R����%I��dL�G䨓۪���2cC͐-���b�/�М��L=�A�o����}����`��z�TQ�nұ����m��TxhR�DP_b�ld��yH�f�)tp��>���E#ߍ��ǌ�pӥ孺D����	���}�c٪�5i������5�K.�rbi���S.�(	��)��ʏ��i���3j_dӵtg����A�+���5+/g��XR����9�Eu�v�H��`� �&�"eÜ���2ܟ"		y���C�UL�<h|��.��5�ς�p�8��%��Eb��]]���yGvk�������W65E��Z��@C��x�uXՌ絘��J��Ķ�k:H�����WJp���d���o
�N)��wG�A�:0Ӕ�q	�k�<oE�8�PS�n�Ȃ� =��^�c:a5F�o�����IRdZ{Kg�!���l�ۋ�w�*��T�<b}u��@�cx�ו������e`,�h"i�	a`�;(��J�:���jE��$����n�<�n(..�QgN�^��_�qKU_TNNď�ؑ����XJGw�D�=��s�	k��q)�������n���F��9>(Ywq�����KK�����v�=���O,w��ma���&($��Pཐ*��t�D�ľ+�8V�oZ���n�ݓ^]��y��q�8B��C���ʶ�ë1�J���@��W�w{�(��|�^�+si��C1����q����\�ӥл�Vj\
��-l�׾>���̸���5�%�G��?��h�Ԏ���5O��4o�(��:	�N2�\N{�A��G�-v��.�ywy��P *I�����L�����+M�U��my������������:Vu��K����D�#�iO��R$�g|�$Pi'��M��63<<#��Ɠ�0	�<~^��?E8Y�<w��2�~t�bP̃:�j��o��>]�@/����~��S�N��P���J�k�)xv���z�>?��.�\c��O��"�����gΠ���
�#��P�N�������&�4�ʉ�B�?���93��a�]�%�u
ݦ�-���χF��ǵ�c��qо�+�Zwň������Ԑa4��O�@lԍ���Q*����y4��_x��Э�;=���׾Z���A!*)���}*@ղ�\L������b�(ik�/����7=mű�S��T@HDTU��X:0�Dx}����9��l���^��J�>����� )�L�+Ƿ�:wr�����Ӄݵ�،��&ip�M�Y�$%��z�1)ƥ ǵ��������3�������;��շ=�Z�w��oy�=HS�V�ֻ�d!%��0���c%��\�R��7X����b�͞.i���)td�P�n_�����@���N�9�C%L��6aj�3P��
q�9��T�����
y��~���>�+��<>Й���p���ϘO�Q�XZwvb��ʝM>T+�fP�߿o�D䙧!Cڠ~��=-��n�y�r�O��.2�� C�*�ƜN7Goo��ǅ=�#�ӣ�����I����k2U�b_eJEF�t�����3SVM8u��;hX�I>�]|�=!B��A.�%-#!a|QRr����_�
"`.!��zt����Ǻf���?�1�y�(�9��^�(>����N�f�d�K�+)���-����ND��:0�
|,wo]��g�~r[���,� �}��h8�p�Jf��Q�-���+WWe�ˠ�A�vL�զ��,�J�u��� ��}�wո���*w���?>��=h����5!�By%H���{�%3��������OdZ"��D G�-BH�-�i[cFM��V��hȡ�;8 �'wF?'ٽ�,h_t�D�,IV=#���;�^H�B�����zs�b�I�3Ow� dE��3��kj)v��0�Z#8�P<Է@�X�XIPq$��R��Ή�8�sR�}�k�c*�6�����ts�"��+�'CyZ�t�t��(X��E���{��ɠ�U턜����ǵs1j��]����nn�S_	�G�g񀘥m�=#--lp��|��Y�n��(�6�=�-�,��xH�ع���T;ji+�u���� -\\��	������TH9:�	[�D &  ���N(h�?�42�{B|9�.JJ�_f3D�4;c)9W���wr�e�y�Z�Y���|򭎯���U#@Xٞ�w�a��z�)��2��V9�F�CfC�#1�����Z�G���g#mH44�����/����g��~ީ���f��������|Fژ������\��"p:�[������K��N{�`��f��@���}���|�[���I��/N&�P;|k�r���,�\��9�b��	���b�7W��;������Ā��w>�j�!? �.�gܨ��G>�b4��㡆��e�s�WRh�|�zն?�MZp�R$a�_��6U��{#kG>�ZvH$Yt�X��p���0A���/#5>��s��<��C�x����}8���p�������Ǹ�r�UH�RL�`��`�@N��3�����^Q
mJ���k*����g�[�Hķ�A@��ܑ��.z��|	��<{.�055��	���{\U�q�n?sb��Y�p��t�0>|��<�� ��dG���S�Y��
1��T�֛�6���jrh�۲��4ҧT�9w�'����;�*Dޢ������L�$��ȸ�$�kp��S!ޓ��5f��x�cr-u%~:����@�@�Ix�@M�\�u�2ի@�o�z��ғQRާ�uK�����Yg./�e+��%M˸�Cw䋮����)4��ʛ��S�l��gTԽ��١�ˀ��/��DLWpZ������ϘؠbX!а�� 4���C	�̞���`T����^Z���qq��L���ꠅ������?�Ro�Z��$z<g���I�9Z�G���4:\�b�
t)Q����"�3��=�������̖w�I��X��> �K�|��E8~���?F	������yJdh;��
_�������^�����fN��O#��{ ��������W_:����n���E��x�>���ˠ�{��MV��I+^-�J��m�6Z��<M��ށ�k�|�2��"����N��ڰ:�#l:�<Iz9x�[VI_x����u�7�o�bt,ʥ�ߠP7}���JJ�:�1HNFv2Z߄��K��������)�%%�15�y^6��^0ۗ�r�W{~��u�O�ࣖͰ�C�F@@>� U���l�gd̅M(Zk'NA8x�,���+�Ag+���RR�5R8�&�Fȓ�LFQ����i �Ϋ,rd�O'�?4wݗ��휡wʎ�����o��g<�G���I�Aֶ�AV�ʉ�@Ĉ��B�d����M��>�:����k3��I6Y��H-o�9�=Ar8��[[<)��8p�������x{�֗���&_���TR����D\A��ý�ۀ߻�x;��w�:���_Y�"Ѐ��)죦�(͢"���&���dH��
�4'Y�Fn4�'%=&���L�w�SU���zxuk��RU��A��7�_�(�1D�0%G�%V��4���
�:/�&R�`�7T�|Ñ/ܙ�l�����Z"��=�H�P�C����PS���ʅ̂�@l�u�l'�F�?����Ύ��;WMm�~����7�V䑙(�������f�,ll���A�
�M��KemoO�S�����3F���e�E��7��2���g��k�c�SH*b���k�dq�p�AS�C�DC��A���|_�6E ږ�{khh�$KJfA������嫠�=:�딀���������P�J>#4��2��v?��RzҤ�$Ǭ��%���!��R��A����a�1�q)���#����*#�B~�1�O%Y�/���}W���z>���Qndf��lBl�=�c�0aɌ~�3ʋd�+��Vp	|�d��1�E��EQ�#����ݑ̐�������g���`�"�d\������{.,�(�Ʀ���!�΄�9��'�@�����f)}�;M|!�ijn���ε�y�bi)İ�5G�wvB��YOt5*�լ,�������2�cE*�yt)��D�_���;�� [�����r܉<z����-H/4C������=�ݨ�r�ڹ��%O$��;фߘ�j�Q6��:p�|�(mB��tyX�[Ф���_�@x���X��_U��vw�`R�m�����0_�4�5i(�£�����?��`�j��ꭙޤ{��,ͧ��˹Is!j���m�|8��n3�Iw��}ĺھ<���O��śĬ�Ak�x#��ۮ�e�9p���v�+:S�\� ��f)Z=~�\3>���/����WKK�����鞒1�3�y�s);�G�uu�S��k(�b��W �ݾ��r*gPl����en[e*�x��>�T����uM��HuUCK,S���;8s��x�wq�!;p�u�%,�"�@��/�ފ������� 6^�dMB#힘&Ĳ7���}�������NJ���P�!�?�}�t3�w�y��Ś�?�fe-�~�al�j;d��v/f�	��i���2�C�P�����kFFС������p������g��0�(�|�@tpb���f�3��n����(��(P��E�D<ˮ�P�9�{G��`��w�''a�koݴ�? '��G"wTe�u$�߸
�ii���G�y<3o�%�K���HNLIq^(w�r;��I��#�d~�
��׻�LӲﴙu�N������K����7O��4�)��}T��� �Ȕy��
��-j�A���!bCF7��no�nz�ה�`�X^Ǯ�Ft��\�Q�Z�?V���Gll�ۓA�EH����X(i&%���WcV����b����;�8Bŀ��F� ���hfU�m��/6�li�C0&�QG�Ë���(()Ü�Tg�]&�`!�� ��$ ��J�(���,L��n�2IN %�O�rp�M�F��@=6�.�=ͳ�[\��x����d�\n.*��(:g�_�!�M[,Mh���$�>�?���0�D����L:S�������@�a���-b<.~=�pff����1qzA�>~��Θ����c)�	+,v���t����~ĸ�q�SS�C��/(�eQ�Aw��	��Բ�g�y|�Y�d��=��[8��u}���97��>k1WPXh]喾���M>%o�J���㒕�M�Ѱ��C*����	�+1�y��H}��kd��o+�"�"6�җ�m�&�|Gp�mk�2k?x���y��������j����:�&MM�zHr!4
�©�e�>fP<��>7���k�;��iďZ�-(|BE������O��A�.���es{���a��_�U_�FSrLnYߠb/1.5�8���6����v�?Њ���aVt'g���
�.��Uo�z��Xw�Iev�RU�����}B3B�����a�be�* k�i�§=�
��v���B�����5UvD�I��.@��u�Ɯ�_���W���w4E���US]v��+t����ܿ�}��A�mȰ�En��Puu���I|�������A����w������GC�H,����rPKqD�0f��bb�芖TϢ#�Y-�\ǔ����o�B�����k��ލ��O���_&�B9j|�+rm�#ǋ�B�M�feл�|(����6�כ��>�Xp���P���\\s��U���)�n����3@6��A	�.�Rj$��6�EI����Z�rn�|a�����A#RN`$n�N��5t�l�m���7X�TE�ƺo�zV����C��&N�h^�Frh�*����樽�G��32X��O"����o������iۉ���r�;�<��J�h!:��u,�MLxI�����wd�����[cu�^��W8��z)Y����Er��=�T.�et@Gm?tG�!�\8fd��rÓ�kHj�-_Q(�G`{�a���7��  ��}�'<��Pp�O��S���^���4�N��� ��5.�����\\o*��Z��������e:�����W�R�����Ç�;�z�w㔄-~�����i���~v;��ú����C�ml�S��F��2q�f�b����HScy���z��]���Ϊ��r��jnO�P�|�YD9�$!$�>>.�םb�C�V}�Z����"��+"%Ek+�B,q��^�^^�qj��n��G��bT����Մ#�C�����G`��s��(od�C&Q#��~��~��� T�k��jb�&H��:��#"�kv5x8���J3ā��fmӔ�J��ZJ�T��~	)G��b�w������������o֣߮�z�w7�e+�~���8�5`�|��\��
����j�h�0��B]�����}z�w�L hZ91�yLI�C����c��b��g����[�u5�[�������<Y��� ד�1�
��LDD4l�<x���}�4`c�l����-N>�����I���'�踴��-s<},��?��r�L~�X��]�]�U�T�8�v�;o�J�*�Ƭ��x����l��e���=�������.7��"�ւZ��j�i�[" .c}��-<f��[&ER�W�H4]W(�.���:�r�����3XT-4�tlE�.�M	��n��ncن�5O��޺իF� ��iZ�Ĺ������ݿ�Ƀ�(��͝�ۿ��#>$|1�^nF]*�k`�ƋXR���y��b�j̔���[�z�|��Q�Yx��;-^P����݇�'�^�Q�����]pR�?��߷n��i��W�������=�r����ǜ���A�{$��Y�6�p�-'U)�\����|��Nt�b2���[���Z[K������
�¢�}i�wJ�W�t��N�a�� ��H�d�Ι����ˋM�L��]8�T��֞��w�V���_κ`Fƻi�)�Z��+C̕��ۀ0��d��!��-.~�p�Q/�gmv�nG��V�IB���&�,��HYA:�uٻ��O���?��ʏ�md��\&H�ƜN)���6j��u���mo�0,���E">ߣ�"-��AG�1�F�fcnF��K������z� u�4-^-�AR��Cy�N��^o [11�q���b?�S=4�<`��e�����_�3t�:W*wn�'���g�R˰ B�Ѣ�/�%?	����B����7�}tG]\�>;<�_�|������:5�y�H_;�. ���"eGX!x6���ȕ*"�u%�	����@Ha\��8��]:3U@w�G��o�z�|+���9֥"�u$	�]~�ʝ�V��w�!�67#7}J�:1�A�L��"W_
��=ٔ�7�{�\�9�'`?��!4���z��t��?_Ҷ���iQqP	@�ٙ�C	�=�fzI��.��B��<�L��[��R���T`�w���(���xRcVU��f\z�z���T�����n��\?]c�S+�sH)�ܰ����Tb�)W_��g����q.A��W.��0.�]qI�E�b懲�u(F��ȗ�CM7��wPr}u����e��G V�)5�}8�����!U ��LLL R�f?q~���=s]?V"��,q��QE�$�O�ax�K�=<҈Jau�� `��p��טG�G�v��z�;Y'k�?C
HjŎl�D�IE3nŋg�6;����=��SH3h-�A�Mդ��%BSU>Ħj�?�0i(���#٫���z�%L����3^
zƿx�IU�I����1�Rv�oA+�)�CZAs�zA�n��6��Ӹk-71s��QiJ9̂z��knV��;T��c��qmU�(�KJJ
+l>G�@g�|����{ﹰDs�+��{\a�o��� �#�@;�T6�\-3��>,n1b�����i�; ��JM� �á#):��e�ML~:y�g���i��
�5f��^��)w6E ��:6/D:u��uȻмoc9)aq7a~N�XY����)�WS�9N���5�2bc#�Ԇ��5A�)?�kG���m�t�e;�θ����d�!��(���s�:���'F1��:x����zo�]6�8�3"MGW��#`3��F]������7�$/������eƤ�e Es�����edd�Û���g�G�G�����''lϦ�"�oo t���!8�"K��b�H�y��T��IPP��P�I�w�.��	��h��ѱ�/�Ņ�+��=;ğ �,x~�C�@5���䤗R����8Pz�S��[���E.�RѴ�������s����ɂ�[U^]����gV�=�!������^o�˟#>'v �{�4��))(>��(G-	⭪z�ܰ�v����n��	7�9Jw7�f���o�9V~'W-��F���*�<uy����!-�+-��c���Gm��+)$���Y�l�V�w��v}���gc]�yA������{{�u>�ƈ��<��:*ѫ�#�J[�������"��DЖ'j��e�+��v�mjw��cɉP��	.4ꥸ��pVK�b<�U'b��S
�P��?;o�k'���OACy�� �Ӫ�o���"�lR~=�~hXj��N!i��a]�q��<t5W?hߏIp�gc�}����*eoo?��؜��Ԯ3��!����wHbk;g���2��5����Ejdd�X��F�c���+�-��Ⱪ"� ,v������� �g��tt��Ș_G7�Ck��qn!��)Q~z���Zn�g�9�ɖ���"s��&�*�?47�Z���{v��9,��X�*�WJV��PR�Vq4�E94�9՜�6�{5&��n_�3��~�LO}Z��O\:���{�g�`�C����P�����6��ه|al3�?�^������I������3�;�)�(()_k^C�4�
��*_��OL<���%·r��=�"	D���#Vټ5O��ʘW�ZW�X	`fUU�P�&4K���i�%�E��S�0��s�P�0��:|�L�KK1�9�L,,��by&Tj1.ė��"�d�/�dx)�/�5`�O�/��w�/F
�C�q�_�|��]�u��]H��DT�;xQ`P��T�%��֭4-��Pg�|�0R�2�#:�%��Ӵ�!���I��@�P�,�<9� ������*�O`����b_'�E�b�v�׳��A���k��px��Wcb��d�#��lWUF�6���������>���t�aZ���@A*#�3�}7t��j@)�)��'i�XIz>S3y������1|9�F������� �Jfx��|	D�����*_�>:���h!�j�ܜ������H_�]��;	hq#?o���j��U�N��ʙ���^~�����m�}���E��^����m�
��*�q|���'�����!�&�4����Ҩ�K@��D��ԄԶ�V��.a.��А�4�&]YY��� �A�����z�/	y�K	=�w�B`\8o8*ιIS�TŠ��h9��I�b`r

���!ó@0��rCS��n�9�[ނ���[��B����wO{DV�f��q�]�5DZ�mO��������?KY�	y}��#�r�p���z�mH �����ԤW��VGˀm��8U�s43颰{�K�<���%Yu2%�6+�)�}�FKt��d4|-S����y�����o����^TZt'�$	�R�R��~����^���INj�,W��I:�k��������J��9www�t��[\�1��I�w���\޴�����
AK�5���΀G%�K��|�]j���'c�܉�׫9�4��1~�2�?�91'/n]�|��ɍ͓�c�"��~�iB�Z*|pMsꚟOFbgf���ř��Hl����ǜ@�zhF�|��O�����~I��]�g��x�|`p��]|d$�ڦ*��2��ݫ��@a&�Z��y�;��a��KF�j===�H�9��"��T���'dn[;A��G��Sw=iVx�""$.ŧ��G�6�q�{� �ԩ����JB��7�*ӳ��z@*|i���7�O���p�E-M\
�[��p����������U�5����_ye��VH��[X{�J����oət����\��\̠J��~���4��Ԥz���t\���Z�T�5Q��`E�\9�I�B�+��)��Pq���
��	�B�y��k����&8���'��_��߿�A�W07��eb��/7��e��R��1�DR^F�Z��Kr����/����i?��5�ξR?�"���P52��?�-���p�����!K�9����|��cH�6�
G��pr�'i��Q-�����s���݄uP��=���������J�*�O����55A1�0�����-Z�(�*pЂ�F�}>�b/7בmaa!^�}�s[�P�R󽳲���1�.UO��m��Gf<pB99I��x�4Q���� ���̀�u9�h'��Q�^��_�NiX"3:�����R겙)�޹R�l,w��/]^4��u��(��Y��i&>�ٱ���T��+�
�=���n���_���u��-��ݣ<"r�:������DԤ��qR��G��ח�f���ۖ��A�"��$b��������C�Q��{�0��r�aQ�����.�^�������M���%�[�hh�ɠH;��UMMןS_�"	#ׄ�.(4���75��Y�7(�צ-gfa�n�w_�}F���
��o����Jv/.���BU?�tZ�`��SDCM�p	�J��#�?��wB�w���L
�<|IuKU�re�枸��8�Gd�ڽ	xR�,�BY&4����Gh���7|��'���z����Y��C;'� �	h�+ ���J�=,���>=vL
���I�h����Es|����axw^�Ź�KEh ��&��""�X���(Ɋ��hi+,L��x>�5+��15�:�H��4���̴eZ�(�K%Իܡ���v{qw ��(���%����xH8}Rx~��b�w$[=���cڹ��8��x���u��e:-29�	�O�D�`.��Gr�F�<���C����v	�a>�ԏ8�ډ[�����m�0�\,q��)w?��Y=}J�P��:ڧ׵��q���Ʊɘ�Ɣe�aj�Dj��-���v�����^���t��%c����2˲-SSc���R�V�R�/q�{{1:#&FR���.���Ѥ�{ۦꝲ#,D��3w�Ծ��§�/��aM��^�鬟K�
�`h!��b��O�́���+�3���C˪9[��s8if��j�f�[�I�^�$��F���NN�ߪ�{`�o������ʱq q�J���{�eDR6.&�Q9J��M`[n0.[Xx\���_>�wH��M�&D�_��7�,��^GF~Ө_PzX;����S���eR"5�st$ ��\[Zbj���/�Ё�v��B+�C�KJ�e���mk�n�˻�������Qq\�_-�k⚰�?&���5i�|.Vd�5c]�=^�P����)�J��?��Kّ��?�r\�d�2��!���κqG��v������w@N����F�©�?��d�Ƭ�N��X���N�Q��a��}x��a=�b����3�G8� $�Z��{���,��o�+�d�jM41]U_���6E8B���X(h���
!�����;��jtu-2��d۷�\.(��Pc6\32r[�]3�H���b]hi�!M\�����&�����y��e8'�W���[�j���Q�6]��Vdƃ�a,�4-�����E�t����Z1�>mr9��Z`|�W��Z=���6��a�ݽ�Vʹ�v�c
^JfXS�Q��G�jk'����'���������k�	!�m�z�G����|�����K4G���@@�-�gfޤ��-�<�Icg��.u�پ:H7KqSJ����	l�ņSS? ��'��y�Ȗ1�ħ�
M���Q�,��AZ�w*Ãc�!.������1W::�	��4�[�ir���5�u�NsH�҆��e�)��߳󭕪ܚN��Q�w&r�=�)���Ż�S.��g3�RvR��7�W����UMlC��R�a	_�޹ YcN��<�:�>>��
����Y�|�I����c��{���C��/��r��l��){�n�������JJ�s@���=�i,���!����wh�WU1pr�yvK�b�l͞(�b4c�9�m,A)񇠤�Sb���=:�����L��_�aۆ���!mxl��Q�,�ٟo�ko7дC�)u��q�uSoD_�\��A�����L�Z��K�G��Ӥ�3��͞8i�{mp�3��!���.����i�FC�߭���GЛ����	SP-̾NL��`�Y[�����S�%γ�i,�P�BLX�Ga�E,�g��<a�;Q��Kz7j�n
����v&�5��>���'r�Jڏ4d�G��;+���������;��Y�0�ͅ�l��.e�� �S4�_��ABs����=�C�$G��j�R��c]��mn��"Ɖ��?ؒ�1k�s���dT�҇��AXFW�w\jU�� �=ʼ.�B�!���)v�3O�wS�R	���4u���!���~�H���F�;�/�-�fҁz:�l�$��eirg�_ɺ�0�黹��E"�1�++�"o�^6)6���q�2�Ihw��K�Z6�o
\��Ov__��Gk>�oA��TP�����q|�"�t9��֖��i^���d�d �
�9?CNFF�ɂ����yf�5�Y2���v�-����
��Qp��%��]���=%K���<$P��"��mP'�}� o[�2'כ�Q<lJ��@�k+�c#U��Q����}����S[��.�9�韭G�B����dZ���{]E{ ƭc]M���2�1����Ɯ){+��$�p��Υ�]sK�g�>M�|��b7�r�Z{6�����,��ޕj�+k0{&�HT�%nS��[dbh�����{5�ܾ]H�|� Hc�		�΀�G
G  R�@�x�3	��o<P��Ⱥ[$�,�A�km�"�8�=�����u
�F��+�f>O�f��_�Τ+Z�E���qY����Z,�mjty�**��2�Xo��o �$i��V�q��4���ͅC����i�#v��@d������M���sjc<��m�TP M�r�2���W}~s�ב>�..l�^�H���nj�$$Q�GT(��,���Q���'�޽[}.��B���r@y�MP�������֡q)�Ck��ԋ߿>�x�s�/�@^������;|����Z�e�~���%���f���tk��i.�z�#�y��g�ܿ��{N�e��*�Y2p$�Q'uom?�lè�h9��l�yDV�v��?-P�W0�o�y�=�g�k�YY��a\�Ω�{T'a��k۷�f��k��������p;�����;��;��7B0�C?ڣy�f^�"\@6P%���<s�)��h�Jp0Ć-��ؙK�l|JI1�[q�QW�x;z����>����a0R���-�~G:��gci�©]h�������� �X82uX���%tt��ϥ�o��7�6�g+nR	0�N��MV���NM�rr�f���2uH���~��w|�4���,h}_l���q��qZU����Cp��U����:~'���yOu��'�qq����y���BxJ�J�
?�XwB�?���]O*֏���ww�"|��3�V$��c��a�Jk1�A�����E������9�G]�]GǇ�jh�g�������$G_~1.�~��y�~�R&SD��m����ƀS's�6�jZ#�a��^�"7�h���a�P=�D�ӛ��??D�϶+�SL�{���d�F��<�o�ڱT��ToI��@3u
sͫ+�N䮑�f��,�Mcޝ��u��C�|��\Q���D����x���� b�f:�RO摢���3/�����ǎ���� Y5uO�Cި�g���c�����j����WUz�ȿ���|�����=z�(� �=[n��i�{�9x���߆\k��-H���r&�*S�ۏ&YL�<Q ��g�@2��`n@��:��fk[�:�xo�[�� �2�@D	�v��DY5�3 � �[b���h\4⏿"�H�Oh�
��V�S��(��σ@u.�8R�E6W�#��lE���Z�<�ԕ6^L�&��[9�zPS]���ƺ�\��)�ᑾ�7�߿ �{>���s��(!5�BjiϠ8�iVAABq��"x.9����n�a�[^î�Ы���\����N�����_"�O�C��$�F����%�myNz�70���J�a���������m<`�'KꖜL�{���r'�fwq�K��=�SIA
�~�5��u%>~4�7;ED�=#qhA�l�G���2Vf�����yP�ŉT~�ٛ��ba�"/¸|~�x�27���������i*)�6ݻpx�_Dd��ߎ;�WZS�H�LEI
 �@u_������*��2z�J��������	zu������Y&��C����L����E,�^��Ϧc���h/t6kd��ODD�r���(�f.�?~֠iĐSM��Q���hypȽ���,i%V��-���E��B�O������?z��J42.���j���i�x��@]>��h[^�r�����Z�q�1���18��0�ԮZfA&��Q���1)eX���*��G��d�UWjN��1'�yv�RW�ć`q���iI�CK�m�|+�X���
4 !vf8-�����m$j��)�f��-Ⱦ>T��}���Q)��[B8_J��4�qy��{�[6@�p8�l�{}���@�uzZZ[cVۚ'��%��֘��̿�����k����CH8ۋ��Z����73o� ]���6��Hj)����Xeq����~N���q�K�<��QFbAE�{�����M.��O>���W���혤����9�A�-x���A�O��$�#X��=�V��;zs8����h������g_�:�)��J��E�yU��<+��e���"_3ss)WJh�M�"����y�!3�%��aSo�
�.�`�{}ccg�T�*]��ڄ%�#;੟H�bG���nK���:1�|�o�3�*�Y�#�|�	���j*�55Qj��徛�A3�2v�Z�q���J�<$�,��Z��ӳĜ�$�:�K��ۇ�Kfeo��W�Pu��1��7K\���d�9��߹���ڗM����������J�:��O���N\�d|����Yk����UP�z^!�F�lsII�L�97�N���֏Q�u�.2&;��ɒ���}�N�8yc!�\��O]���%d��q8{ߏ��K0� ��Ͷ6��&�>�����W76�_�/vw+|�x�Μ��A�DW_�H�ΨN!iG�z�9
51����Qg.LZ���������˱tM�G��J�[8~j��N�*S�}�<��≵�!�؆�*F��u���x��	D�2�B#�������^2��]���h����?7ܤ�-I�8/�{D<�4�������^��F��%p��x͈{;����[|��	?M��T�����v+��������=����P�L���oxXl}*�E-·��Ts7��0(�)?y���t��rr~�c���&��3�]\�i�aw�}*/O���7N&��_�� ��X��jl��3U������d�v�a�g��������c��rܷ���%��h����bB�I}�>�0y��r��!s�/��WnG>G����|��x�G�?y�h��Z�}uHH/���������~7��{�M���kb+ѻD�ND�-D����G��-�[�&�FD�D�[��}�s�8�e<c<�^�Zs^�k��ֺM��$W�PM[���������[g4 ������kt�6�9�����cOψ�h�h�\��@'�)tR�X�if�7X2,N�+p�c��� Y^C��Wޓ��i�^)H�[Ě��	x���ѡ��(9��(�7�74pm�\���n�R�$�~������Iz�|���_�����X:
!qJ�J��,֏��2V����Pm̘k۸!f�Y���̾��!��I�L W�Ұ�S��b��I�Ќ���dM��{�:=������`�k�X�Ew,';�Qx��
��@��W�KH`��D#�d;��#L��C�Q��s;�󬽋��gZ�z�3n�8�3I�;�1;�mW>?��R�^��$�"i��pK���t��QSW����J�����q"�6+*<Z'l��`e���0���q���\��ҙ�T���G&�(ǒ[RUђ(�Ճ&ߔX��U�� -��iN�\ނ���S��b�੼`��SD�c�*"G��R�c�T�h�ݦד�ԒI&~����nlz�y���G�t���h�xң���*ݘǔb���tGg]�������#����o�v��7ˡsT�e�sM+ӌ�����ҧa��{w�'�N�bï�I6���i1��c���/�F��N~=���Kx8�?A�T �����l�������ߗ�`�+�~����;���[y�+���g��"ECz2��/��������)1�SY䐺�o~��O�}��פ�xd�z�������=̽9~����A����:��ݝ���L.o�9i�O�vk�u.�8�xB��1�R��8@���ˌ[M�J?W%:�6@7�MM��*/��:�5�7�-Gj��9({s;�'����݄;֙������M��4�i�i+�hiU���-���X�'IQ3j�HQ�i�c���:�[c/���7� Ij�c���L+0�ؐ.�0v��T3��]x������s�Qӓ����^+�Sh��s6gf�Dn�N���,�]xe�Dal<�rtûYLra�� ���K�}��`x��<�����gP��F�jλ�m�{��AKX���P�{Ѧ�
��GV0i.m���Ğm4��6��f5 s��Zl���][�O����8����ո����� 
7�;:�:��s�tv�y��of��uv�*�Sz7.�#�:C�,�u.�<oSsQE��� ����LK6GD,K�ᐓ��:�;��R6g����\����5�z�.�/�~^9mv}ƙ��ӥ�T�@����t���Cf�A�â�����6*[���mEYs󏉷oΆ����}�l6���K��5�]k�O]b�?{����oZ�q�2p�	������T��h���'�j�v^�O��2xJd���@����47�U<~2i~�C���F�lU��J��Q{�VI�u~�FSk��t�t�uG�=)�����d��X�O3H:�݄�/Da�
���� R�D5��8Gt�H�Я���\9����-��L�L����;��}!��  sQ�oJ��=up���%��2�����w� ���T�؊ê�v;��9��~��������2���=����h�`���)Ѐ��k�vt\|<Q9ɫ�;/X�xn��xkr7�G��w�I3yJ�N	K�n�
N(L��q4OM���Sl���Č��[D��� �CN�!~fi��֚4ɞ����A�AΛ�Ɗ2���c��K<�
�XJ("��v�g�t�i�f�7c4y��$U�{�/fc�S��#T�W� �g�=֋m�10pG2��_ں���NM�$���%���D�n�w4�8������QJ��ȵ�c���B��|4PȷX�|�& ԡ� #���3�9u�����?Db��_��~&� �r���I*Y�ʊ��9W#���E��n���S�Rn'��N�k�f�����P��v������$_�W�D/���0�8[�x���c5�59�Td��Ԇ��anT�v����?���ha��s�zn,z��D��x��S(ӋFP����jUlf�|�###�����>Ûvu���y�v��ؚi�-�h*?���*fi>7�V��m8����a���;�[�%bP�Ҹ��W__�R �8���p����$�}#������*�4UD�L��`Y� �B�s��M�"����[�q�KȰ��As��bX��N�EG����K�Y(p?�����۲�ɂR)�, ;"���T|D�]�?Bp�V��U�EI	7�����?�@������/��ݓ��񕑕%̶x��񫑒vY))�� m���yx�vɓ��z��쑹�t���M )�]���/fFFK��R��I�����F|��E���~s�aċP�b��~EZjꗓ��
�����=���]�)g�o�ɉ	n	F/|�r� z���o+[gm���1M�cR�׼���w�&����F�}c��!���{��+,b���e��hN�ui�B!G����F�Cz�<�C�J@��D�2��>(����h����$'�Dm@�paa�=Y�Jc�	r�O	―~����1p��C��b0KVỈw��y^��������m�[�����Q�S�o��_]�Q`5�I��r6�:�ƗL���M��3�CJ�W$������?�r��1�G�<%��lu�q榕������sˮ&!��s� ���h ��ö�N0)_�$e}5h�G��dN���X;n>.p���]����41���׵��CJ�vE���///O���q�& ��Z4�a�n0����~�@@�����G;�=]�;�>i�B� �s�������N��_NL�Ȱ��P|�*G�o���*-�x'CF^&�-������f�b����/�bwd�wvh�<2��-��rۿ�Zߊ83H0���<�9�`��0���І�~=��wvt�֗N�s�$��Ls;l1�7|������#�T{X��5�ʓ��i6�D�H���5	�M��ޅ�����`��KX�jq�u@�+���P�O6$%(i:��n	8|����ǜ+f�v�u׆�䤘����nm�n���z�#���~����
��+n����䎊�''��ι�{y�F���9�&�]X�v�W
�0 ?b�(�
���`A�W#Uo3*�ڪ:�DSK4�J{&�sx������wu���k$��ro��h��w��z���	H��:�ߗz,�� �$6��H<�>ʴ����r��!&�Ud�%���Q0�oo��آZPa���C�1�`r򉘌��-�p�q���l���ߗE~o�|�<�Ё4ޣݗRCSs�I$���o�|�3��V�XV�wK�4�j(e���u���H&��Y�n��}7퐊�.�R�#�}c�v^!:�8}����8�&�e4Ի�o�m�U��B��-T�"Uoc��(�LIM}�N�]a��[*���fff���)
p�nˑ��I*
R�s#��$LR/
K�_��,�� ����� �)�c�QC#N�"
,��"�S]s�3����Xݒ�nnx̴_�'_D-K�����ˌ��2?�6*�?k�h,$*:W���߽0`�C�mF����G�9�]�pg��A���۫������j�G�s��B��Nea��r��%��M��D>޷
t�FmH�c�ٱ�{ˌ� ���T�v���У����cct �������L[s����s�Ƅ��yU�{&�]|]
�]�����@�K8��1\�oW�`.��������lL�b�W��g�M�
��hL>c#G�r��{'�JJ��h���7u=�o�\��x�,���/XD����=�#��˳&���M7*ߥXMx�HC�"�g�T��ERcF����|���w���T���U��夘e*���R��a��C��]ϦnB�	'�y�4�_Ic���K�x�4b�/95�'w�-ڀmLΑ����&1X�j`�#>���ޜ~�ez�K}��%�B�b��ȵ��(��^�(�_�'�ݹS��������B��`T:@{	�g��Z�0R�im�C��sg
��c������` ���@����#O���m�(.(����|�nEz��*�6f�/�v�~��~���������M�Q�����KV�;+*�x20�?�&0��Iʗ=X�n�j�罯��,���Ƌ��1՘R)�ć��>��ݳR"溔��(���R�O4>��2�Kd��~c��a#�fUX͊�?'�ޡ9܁daN��r2a��4���C�� �{ﮩ}.���v�9~G���?�;"�+-�S�C�Qp��,��C����o��k(2��ܸ��}�]x������cMr�?��l�G�?VZl0��ueD]S��\��e�փ�P���W�O;/5Wd#����7..��IH��eE����>�ԕ��nN7��+x>�|�{|o����h�ܵ���w�ܡֳtY٧k��s8;{�W��H��԰"�r�{��+1�B<D"Fi�?�*�:z{���m�}�-|0բ��ՑZW�\�%�m\&�ø
D*�4��kN����G��i�=�f-�:5�$ҳS�S���y/�B�9���c) |�bꂕw��/߿���8�:
��XQ�\V��MHȓ{`�������S�����ݫ����C+)���&t���u/���M�UKo�Ͽ�����(��~l�ٮz7�n�����ѳ�f;&{�+Ū���9�(�okk�5�1���VEߋ�^���z7�Y�8[���3��140j�G4d	P��^��w��XG������S5�����EҨ�1�$_cF�d����?Ժ6���{�Ux7|å��^�5`����X����[�ty�4��݄���_Ye����J�.?���,z��h m%����%1qq2�t;��¢9�]��55���"��b�?~�4�6$�b�^�����rQ�~_~#3)A?�r�Vf��2	/t�֗���M�놡�YX�4z�X��RT�	HcTrXD�o����p>�t'zIN�wǗ����`�PlZ��@)$�3ٹw� *���O�	�nl����������\m��^����rj}dXD���Ѷ �x{pfs�$�[$i���ݱm��O�Ē��ɔ�����Q�m���'�,��Ճ�����x	ʣ�?JP�y�|wЀ��yڽ5({��q0(��r�ǀ��H�hH�PkC��1�=+���ߋ����[8[ϱ�ttH��#E)�0�G|��= �,W���y����=���}���~Q������*�r�֒$��Zq8�Q�H�\L��e�l���8�"$�5�ހ�������f"�����:�o�1',�I|������n���O�%�_+�3�Q����;G�������
!A��d�>��74"O=<���y���ku�'p%�/{JDQ�_NS��8�7_��h�=1y�@�q�w�Z�� �Y>�g�s9��%`�Y���<mYW��P�/Y����T���ҽT�5��
��~�G	A��8��߅_=�4q���]�ϧor���i0�[LU)x1�{��S33���jf��^�6��مȈ�uG���C�/+#K�z5�Տ��K��v�Q����-���������vՕ�R���GU`��ݗ����>�vc1Ak�)o�'�58�I��ͤt]�c{܇��!��4�.H%r'���G�@2����[��o�����۳��
��Y�Y�$��kbt��R��{q� $SU���m���mւ�rr�o�%%p�o���^Xu��4�����z!��[��-��-:%��2���:��=�+�{�h_���B�3��%m� "66�~�\=3���s$�Cb�O7��l�SA�~�׳[����oI�Q�JF?^�Y�����"�6M�\���L��省���y����j��j�d)! ���O}��j�沆������cuEʉ���"�5��|�[�Tnk i?���k��^��o�ς���[&�vg[q��Hh��#�k���MiR4#C�i�-2�EW���	��@w�<�J�h����\%��s�$L[����[y�BO4���u�ws���3���U���@j=�����S�Q�/�223#���&z�y���XH1/I)(�q�»B���#��������ZL+�C�|�)4`f���')�R'���XG>�ծ'p8X��֎|���_z�M�H��}� ��뇕�=�i�T�Y�8V=%�(��g��ZEt�C����ͤa�:�S�G`a\V���pK1/4/O>��8u�W�;ZW�{Pt6�F��}0~7�¦mgxuF��k����+���I�8�NNq��Oc�����eC����n�z��?{��x �\%��z�
�J��ٔ�	�]�*�����`�i�,�dƧ���ؒ��f�ݮ��b���|�#�"�B�1�0���S|D��:Q+&�p�K��J�v�}����Nʫ���/�6�.��pz�ϝL V���{��cw�fׯm�۲ӼO�W�qk�uqm�C#�휭����P����`��-鬟�������+<��8
�����JJf�-U�0���<Pd �&F�}��mr�����D	�~��f8n9������1�V'�n�W�i��UZ�!6��K<s �d(v󎌈�>��YX���u7�P��^6�@�^�>$�B��b�H \�����CCP�!u��E��,�kk��YV;�|�:(TT�	�:��íYaM���'zt�--����q�zh��SB��'�ij�U�?;�׷�+�
��Dh �xJ�-����	r�4��+I�3*�A5|��!��5aDR�H�����~r K2������9����Y���k���XŐӁF �f9|�č��Rvl�e�0/hB�����ID����a�ũ���	Z���S��Sx�V�-62���2�� '�=�4y؏��H�T��_�3�p.�B����4t�z�V���.3��O�]�����Z�I�Ν�¦�4�w��D�B�w$4��'(��j�"�5=�K7�^��$��9���ǾvW�w��ty��E�(U��JGĬx7;1�B����5K��؁����G�`�g��@.�ly"�yJCc�\�yfFoa���|�nD��/�.�F.GQ�&+~�P�:�X��|���j�Wpp���Ы.2$\{1��(9L/U��3.����W��O�+X#��B�*D��S������x&�ge-��n�<5��ǋ�>Zƴ4��Y��L��0��i3�)P���5D�^B��@Ϣ=�Gf�l,�|�.�VbB"*��^�vͅ]~S��?���2��@�f�оѿ{$�e�߇�BC?��k�|�y��[������^�4����Z�0�W�&-Q~_K�U�K���Gcﯛ��M� ��D�4��qr�7�\�^��O���@(��H��쬼D��}�+�$�srq���h)Ҝ�;S�^�,r*�8ON�Ґ���"���{�ѵ�7߬�A%��-#�������\{k����Ɋa� ��`�3ӌ��8��~ro[Ú���bZݣ�����6�>�FYޝ�>�RT{j����Wȁ��!�'� r?��v%�$r���L��F��*�m�z!Q�����7���������(�)��V#.J+oo��B���ӧ#�Q��W�%�ۺ�?�>�����ke�F\||�_���֐�ŚlAK���Hd�Z!oi,"kPX�k�O�������F�
��n�@b���=���J�SĪ�ȭ�����D8���g��(F
9��[�v0}�&�����mё����G?��*Ddk4��(e���3�Hd�f�w�9<�m�PX� U>�;a��Y��ΐL�@6z�H/A���$��K��B�Y/'��W�b�=��R��mR���M����V��Q�ּ�?����0��;��ڧ���~�7�aig�d\_�OC��W��ŗ����n	��Gc���X�����(5~�D�b~&X$65��FWN;�阱|j������QP��f��vr6�/�{�Y e�2g�}Nh���c��G1������z��m���u��4��«��e��z;7N|~������ U�mF��4���Q読��j�A���3J~��t�u� ����(���o/":��#N���
E�T	dNxP����WRP�GO_���MW���{m��X
p��U�O���tq���ɡ}�7�/X�J1A�#�������s�ef��I7�F�u�&þ�c2�sw��������:5���:���O>�(%���Cc�SdF�������Y�D���1ǺR@}#�����JJ����@���d���[M�^(�Sfo?��ini��O�͝\D@EPh;��]��[�_J�Y���\��'O҆��N��q�a���D������u�ua�K�� #�Ao��| ����l�	x�]�W䙶02����Ä�z�-i�F>%6��"�y>r�3�v���(;t��?k~|#�V�5��H��L��8u\_6pR�^9ZU��	؛�,�J��sQ��� [���>Lѩ�&,6����&ѵ�����u�ۦI��l�P}�	Ѱ�M����*eY�nxߪ4�kV�ٚ	B�	 ez���@%��$:����D7��t�nnH+�܈:u�5?j�ĸb���N� �ؓ�?h&!Ē+�7e���B�ofvU�!)� ���f�'q��v�y����PoZ����E��޷� ������ö`�Rt.�q��a����?��8�����|t��|g�g�f^���3Ms�$H�<����D	Q~�=ܼ�C���
m֍�y�e��4��@�)��=��-),�ظ���b�@�B:�cR��w��G!#+��������4O;IX�u2h�_��%�ܖr����=��OMJ��7�y�ɋ�J���Ò��v��6����4ޞ�FA�<s�*;þ/����>���k�R@��p2����'wN�lLC��])Z�`�F4�?wd�^�90� u����m��>�#{�4E#k����&��֗����ﰰ �_�pU)��77#֦�E3e���ð���ŉ	r4�_�z	Ҵ����pd�M��5o����M@��ܱ��(ƨ��H�_T䢬���~�/�/�Ș�2ܔ]k�9���J��-kW���Û�T��rE��>o��J�q��� ���L�UkAj�xziY��I�q�q��vG#��lm��%hy��s5�d�}ҭ����o l����%&Z��0�E���xfvV��*lA�#��Q��`:�	y�e�h��U>�����V mTP�$w�E��-�rj@�Z�(�O�;�Id���֯8d*�ӱ�[TK�waU�_|C��G�]�����1�0)F�J�;��&�c��]�ȑ}��Mr��J2*��d��c����h��"�,2fc\�P���'��<����#����R���&+\��桻dm��kS)�J�����O�s��@��JV�o��>�D/8�������ml���{s����^�p��eD��9�W�u?u��f�tÛ�<�?p�<��y�81����*7�k���rȠ���x���f�3���]�kH���,�r��XJt	��	����������A�e���ɴ�B���Psv!�N�	�DOg=��g�̏�����䒃T�J�f��������x��g��U]��E(��o0�D<q���GF(�F"���2||�Q�r�O� J�D�g���$%{�j9��0�l�c�\Ůէ	`Aً�O9a�YK�.�*7!�KD#�����&��e�3h�إ��r".̾[��EQaa7�w����	6
��K[�At��e�����i�=?Xɚt��᝚�W���ec��ϣ������A/��HJJ�Tļ�޸��"d��=��߁;PO?�I��P��,js-��I��AX�Է�s�.��KJ����oƿ��wz����	��%i̾�� C_��hr%(�w��/��4�EE��@A��&�:𷸟����P�k_�t�2�I6�&�۲#���9$+{6!#�;W�󕡭�<T�'X�hX����H5	�$�dL�}�8�F�����q�k�|�:��S��j�h�_hQ�gӻ���@��~${t��������\ah+�`�U�������;��5O	1�q����k�?�D~i�V�}_|K���߇e�|i���XevKmaG�܆�vב���<��GG�}}�I�R6&i���ڶ���:�y`����@�A�@g)2��lo��2W��qUm�X�o2�b�h��.ہ�R��>G���
���#�~��}R$K6�am@sc>�*Ж�OM��7��(�I&7T����X]-=2�	KQ���쥆n�GZ�q$v��$4�1ęu��R^��G�c ���sB3�{Cպ�n1	�X��N�}�%��L.�q>��b����N0�����lY��ɨ����e�^G|����c��E�n_(��aUb_�"�R=	����fc�O�f��34�FmHc[]ň���QKMyz:>.9�=���8�>|Q�P�7��U{�-}gb�{��nM[񊹻�K|{<Y���#�����oT�q�MO3�S؂�J��$`�����]19>R�c��`�L}����,�`�'�/�#+��G����^4>mfDf�5�.g���Œ"h]E�l�OE����f�5aqP$,�j �6úc����S�Y:6)������<I�o�;9:����4�!�WC8�f���?/i�ˤwG�Y��Tq�/`0�s�=_)߳����i煱2��oi�s�@���G<e�	|Y����}�r��`��MWW���z	�ck^n*+SSR�|�
T���Ǎ'/4x��^����O�t~�|V�q���ɞ�q+9�*�a����Gl�������!��=�fW����@�c)y9n�N�u/�0@� �G7�|��m������QǺ�k�Ƽ���B)� ���Lѫ��Xc_�g�0��fY��|)�&��w���3;v�p�*�p�^m!�,��J�]o:�����Xw�l/�Ј��� �y�>�N�ƕuk�%�S8MAs��{�Yf�WNBП��������KSb��^���M��MO�Ɂ��ŝ}�?�����H5G���$+:ÿ��P6���Dr�2z��ѐBw0���A(a�\ ��V��c]*���/��:	�b:%��t$�s�x둝����\�;�U��G���߁��y�������!�'7�\��fh#Q[��ve��j�!ܦc�h�ʲG��D��	�����)]I»\��������`��ә��nړY߾ 0�96i����I�R���tE ҥ�� 4T�a[�+XR� �(IѲ��㣵����8����"�e��C-��5���e3l�k�Muj4�����cy97tcek�I4O.3ytOէO�w(	�$$>]y��91IIa������P��tшA�c##jNb�+c	�ˀV]���|��^�S"�� y�`=S�z�w�_�٩��</u�B�)�K�2K=��'n0���:�:��.8��"�΃���f:�j@n���?P�L��H�����C[[�w�<24��'�D��2��xY׮&�xD"ɝ�%�;67~A�̠%�=��y�8���I��Iu764tLֻ�B}��Ы�A3���@�,��pȊ��Y��DƣǏ�
Y��m��댾_��Yɦ��r�^g!��T����265�Ao[���4�iD.�t�O�(P������C�RN��#�~�Z����4�$�P�o�V"���m�"`rg÷bw��1��!�-u:Z͵��#�/#1��{f������I/0���5�qm|u�K&��_�� ���?�E�����A�.�Zk��ң�#�`�)�YC�6����5�>4����x����,66��"�B*�Ĥ��+"��Oq����t����t�%���7� "	a�MEZ���!���T�5)$���=��10��z���Nߥ�����tm�֪����p�Yォ(_����^v�ڄh��ީ�:�EІw���pQ�������*>�|�߶ߍ��FT���5X<���H�`���J�k����?:~ed<��Y�%��?0�3ߤ��rlL�0�yt���������] �?j�|[�w&6I�,Щ�g�O�dH���0�)O�)>��0�����g��8p5DRC������3�:x�h�/p����aqnBC?� �ߊ�/z��~ YJ��J�����:��u�#"���<�.K�(��cZMI�Lc�ZN\[AT嵭����
,C��<=��c�{��xn&9o.7u�2BY���\4�����?_`#�ɑH�cBa�^QwZ��3[r?:_��*�1�<��f�7g�}�k`YRn�����{lB�1�m�.�w�L��l�h��9�V�@���
[�a����lƸ�����G؛��楒�]\2���4�4H���-%��_�񃢑���"riO�bJ}޻9��S`�<�ώӞyy�$����A	�i��=%v�v(�S����]f�ꊡ�2�޳gϢX%���t����*�\\����p5-X���s���^`P�,}T��fZ�)�x��������qz�x�5pS��|��1��������� %C�	: ^�v9������=��l2��--�2����칛�y����C��Q~\}���ǚ�9<����t���������q����h�>������1|��
���^� *x�T���D+�M��^ sO����������(���j��k��{JM��@] �d������ma���XX�;�;������A�]��r ,�oơ�(��T�?��`7�+6������1A'Z	�M�G&��2!��{û�K�^M��u�v7%�+�gk�����]�ul�z=��Mz�R�v�<Ffzu5�w���>̴�N[��D*�c}=����%yk *gs
��\_w�^#�����Au�io7fNN��K2Y$��"���PM��k� נK���N�+�	�-��M>dުC�tDP&��餫�¨=B��ˣD�Ք��'���>��ݓP��P�]�]��Cm��kfC$Wm��c���(�q�z�o"�ڍ�<������l��Au� �aSkJ�Xaaủ�cyc+#ǁ�;[�e��h0Y:���Ι��d�7����"ꊇ��)�[�R<��3��ܙ��\�:����o�r6�A���n�����}�t<��'���
�hܮ��������g+P��x�5/ҚL����,�s��cwH7/�Ytd��0T`oH�b�|^�4O�\�N%�J��<���G{�\Z�6sMU��6n+����N"VPK�l{v���ɶN*�_1^.��(+J&)�kɪ����;�������n�qA9�p��]E�Ũ����⏬��}4�R����wa!!����5��@�h��E��z�A�E�3wnj4���L�Q�b�?��ገP#��D�g���w?v���y+BR������uT���Ń�X%_,��������3�v��?����h�N���Ŷ��1���p7/���NP�B���5�#�WQN��D��ߜ���2�B��y-�����'zT&h{ěۤ�r�N�-k4����y�[� � 1~�/�7ʾPc㪴}��"H��R��A^Us��.G"�^ ��=�:#�	��uV�Þ�2�T~�t��簳,�0�d��uLE�F�F�[���wI�(�(�����r��� �F�u��he:k��8�O25/!KN3�{�n���>2K�g���|ӿS-������1�^��6wת^�M��>�O�^k��,=��i��Ͼ��}?�H�@�~����GxW�����2�hr#{�1�)���^I�<Ylm���fXN!&��"�����Τx�=u�%.�9�k�Q����Qd���C���F�r�����Ų��>Ǌ�[�e2�����D��]s�,I��W~��Hw��7�����)$@�0�)�TF�����[
!�}���F�N	���R����tO���waŶ��"I�:Pu6�w���p���>��l8+��M�*�+=+9�i~-����;��Bf^2�a�%������V���iNS�9�i��ޞ����Z�x�"�IKQ�e��M�͆���1�ԮEnb�yЩU3x����HZ�ظ�,�n�d�FE��E�v�V��IC��T ����l���O}��7���Z�N�x��W��8�k{v!�<_8����wP)�C;��BT�P�Z-���ocǵ�ܓ3NJ�=��7�p��D��V~�,	���w,Z�����{0/�O낱|��������<{6G��	&��(f�������6�C�ze��H�%�FR"< ������A[��b���U��7���j�y�����ꌨ���n�z�!E;~�/)�e�������|��y���,��ȭ��$~k��w���h������zM�H�^�H\yH�gU�UX8J�i�:�lH�do�r����/�F�.��s�_�wͿ��7��:�v�c��i�4�O�#��~�?���](%~:���#t�w��;��]܄�K���#/�4.ѿ��Fq#U�[W8�����5Qq�}��M/'�1t�l����g�wN�#����vv�3�"Vӓ���/+F7㙤�I��x�����K�[9�����,>B������3�3m��f��;����W��:{� OV��k�z�O��Z�j���� 0QK�I�#�+&��όX2����70x��YnҸ�J0Yz���қ�a4�C[�.�;*��'�A"de8(2 �($�nOk h�'���t�P:�����₠/FO�M��s���)��6����eNsN���H�+����t �Un�{���4��[�u�o � <�����Կr�/ٰ"%#��ޏk�`Mo��ӀO�Bwq�,�����"�s�-ػ��赜�MA�J&�d	I`8�X��ӗ�1��5�p6}�0t�`�ÎO�7R�#}�(����K�(Ⱦ��
ߴut$���'�,�FWXD���e{��}�v ��ᆔ�L�@�����B\l\�����֡����q}}}u��hccc�'����˽}}Y<I�s;��p*���8��,�%R�D-�;� ��i>�5��@��Nwx:��J��772�����B�xS[�����$�3��_H�t�&p�y?��Rґ��qo��~m4�y��#}̨@�S��PB�]dn�q6���)��� ���x�iF���<#�C���2�_��W�'���2�����W�t�ᓌ��LNN��>���b��[��YjF��-�V���զ��t��k��i�s�*�6�r���Śbz@oN��
8�T@k&��d�j��XN8GwB.�>-���umb
;
�,�:bSJ}�֡=�;�+��0�Ww�T%�*ec���}�!���Df���[���/�3R��9���W�vu�:����ۋ@�N#Z�fڂ�4<�q֔����|��*�QP`5	���Ҿl&H�ΐѕ�J��Z��'x��]'��(0��Ug)�A�=�n%����D_!+������0-U���N�E��,̥��L{s�?�9����tm89e�Z��5!%�,!�<�dl��b�X������u��^ǳV��w����X��c�'j5X쫙�����?^;C��䣷�W�x�o-����(_JA�f�����a�`Rؘ����ޖa�־�!�X��:�`���R�*�jEB��5�I�6"��n�x���7g�,CB��&��*��X��##���+82��MI����`F�'���nQK�,G�z8q���D��7t�-�v����űc���}�(�7n��R�#���o`�>imj?�����y�d��T�̵�~��y�J��g%z��^��J S�C^�9Z�~$��"��2�1w`te,��Q�Va�3�a�x�3X%��}r2iU#{��&��>$�C�cza�����ǁ��7��
jV��S�X)	�lY���;�K��
ᔕ����s���p~I��X��mk�vP��20@�������P3u�?���.nQ ��I��Hcy&��	:;"2���փX��ӧ�u���r,-��r�\��cS Y9�"����1��J��7�'7��������Ve]۶q*jB�@�|��*ҋ�r#����%h���\2���� 2Z�ɵDi׿@'��Q��¹�lYkW]3�c�����'w�Ѩ5/�Ҿ���G>U��;�J<�^��RcKӗM&��Д�Ԃv��>�/kJ��eΤD{M9�&�~,/!�T����/��`4q�p]��R��o��J���gn:�:D�(�=����C���&Ly�Id�����^��O��$�f�hL��}k��=W�,)\�	lT �db�%Qw�{\�|�=�s"�4����Q=?z3��Dz ��GC�6���K9k�6d���wH�c>��$ߒ>s@�OMA	�^�h䫮&#Ŗ�����~/i5
������W8G���pI5�����<E�i-"ݶ6Ҡ��E�wˮDV�Û�ßX�p?��K�4���]�5��-F~�mF��G#5<�ڂ��b�#)���-s� ��Y���o:���5�J��iSG�b	��D�u�Hd�`�#c�bz��޴*����Y掩)�E�:��A�pF	O����L���==�P�!�����$@R�L���TdUӟ��L�f�H�ݞ�ꩍt�^��(C�p�;�W�`
�Q ��3�C�U@���[��tK��'�n���&j��sGDH�ކ]�v����p��N�$�;�Ǚ�\_7��N��&40�S�R�Ew��-�`�^8�|�~�Att�H�����r���ǖ�-��-5����iz�e7����JY�r0=?{�#	�EU|�=����H��wz�MC�m�a����!��v��3ц'�v�M$�R#�<I��M�	߬>^v+wqt���������/�|��XX�.JS�e���@ݱ ����hAV̻T�P�l��.q:,|TY�����ܕE�N����)R���{�=��5�W%�n?�)QZ�����}��m�'�NQVv����ݦ�蕍XE��\	���<��k;m��4� ��]YbɄ�盽B��l1a���J�R�E����dx�[�i���%B��V�)��G���ל�.�g~�e9�xIH_��}��d�__�"v�Fu�#�X8��q��w\LU�����G��1Ҙd�\��F_@p%Y��x���k(��Qy�8kr��	�)��7S[݉7�]aʟ$2���P�5���Pu��T���?""�ұ�U�8٣8�3#9��(�H������22BV6�J��3�w����?~�[�ԍӹ���|<��u]�Wγ�ַ�<ob'�vF+� �m�<�k���R��@ʝ�:����"\Cګs�7r�X���*C.6�fN�� y��l}�:�IO�S�2o����R��F!��ռ��Q@F⊐�u9#��F���hV�h.�K
0Y����V�)�V5�_����%��O��3t͏t��q<ڪY=��c�#��-��gX1���V��w��P��2�����+Ȼ�z�	�>벢��z�����[��I�3��{@{څF��\�(�I���y����VYuh�����8��l����J�Zg+^��_X�1��_= �
2~�D��b�A|�̢�[�յv�$)�ӬXOㆉx<w��e��)�4+��e������W���uiV���[&u���Ra�=,{(���'jl�Qe���kn� �������%ý�%�t�ЙtޘC�ﰹ�z�,#ic�73�u*��e�-Йtv�!ǝ�q]8I��L�F��v�ߑ��y��C�E�����6�P����4�Y��W����)",��L��t�Y?��[!�$����y�s�8��Wj�]���6�њ���RKU6zѫ.e�)}�M���ڕs��X��/�;}� V������m�߿�KN�=緍Cb/�fЍ�D�_I}x��K��J�i�y���tŘ�dt����)�S�*f�G�-܄���P�^+�u�o ��;��X�$������#W�-�$�����͹�\���;.���ƺV��٬����z�/����"��4*����$լ[n�X��h����Ak��F�?KV�!�q'1���P�+��*C�"��r�6�����2Z�� {�cc��s!V�OB?h�1��I/�#��}d3�/g�`3��N�-��;ԏ�N.��E��a �$k�t���R>���Y��1�2}X�W��z�&A���ѯ������tҴsmOr�fi+V�^�B"r���ik�ZHɩ]*���;#�~�GS`�swY-;mHd���L��d���n5�Z��=[[(벛y�>,,�X%]��q����[y����irE���ٽc���9��hJ¿ou��b�Ƴ�m�c�
��z.V$��~�D���Q�(�F+��y\
H�X3����{0��p�Ha�snW���h7���	G��Ɍ�0hJ!
j{��_}D���f�<��f
�V�s�E�<��u/^�3��o����:u�}�����U��ޑߏ��t-�+�=�'�ҿ������d;-����n�9:�yR�뗗��Dk�+�ѧ�+$#���D$�j�Я)7���dYu��nq����W�A�VF�-+���cP/���9;\�S%j���|���&�Y�?�X�O3a���'ߗ�I�057o����6e����}�n�JnM�� ZG�	T�/�Ɍx�F�3�4�fOڀq�(n���#�5<��$�F�k��~��+iLV�W�����V\;�)K{:;-����z� ���`��QF��u��3 ������ɝ�o�$����t���d�'hTX��nI���δ��� ���]�����GT���O7���M���5�|3����; ��<)�S��{���u�2��nթ�l	�����s��|��&��T��;����j���L����ҫ/�2���	�ͭ&R �����+#��x�e����ڢK0͊�b����T��h�K+PI��S�4�׀|�)���"�m/1�H�`��%�>�_�㭮hg�I��klW��I�ۅ`��@�S�ݢC8��N�o���m���L�?�������{!�Ҁ�z����\\:	�q��f%��ȶr���]CP�.���!�0	��&$\6�k� �7up$J�׉��Y�����'�`.�����gS��%�'��2��?�D��N�Y?���H���?;?������m/��G�)��X�ʱϏn��]�b�|)�}��~��E��v٤����c���+��F%#����i����ۮ�!�I<�h���5N\vְ�>D�P�z_���B8%�eM�;�����r2Q=6�0��}	+8x��QGl�`u���NB�͗�	>&˘��A~ͱ��Ԟ���y�X��e�]i�jo�G�[*��-π�a�������4tZ̪��R�-^�����̩y��G���M�B���ʂ�Z}aa�l�w����e�n����'��J�C���H$�TAg^�]�~��5@w���H������w�sN�/�L��"ږ��iپ��z�7����3��^i���H�2�.��aD�t��#�ҟ"��k�4}�E㕡��7PI�
5f�H�G���!�W�/��Hר`g,�������hX�=*������V�hc)�F��_�grgU-����&k�1�{�	$iؽ��3�0i/W/`���r�C�4���A���&� �0���V��3ir۬|�@����Is\o��T���3�6�$�'��rzl�X��8u|��߰��NE}�
�n���2wK�Jt@�+�3\���쯨��IL��w���N�c�O�G����G��Ľ!W����cͭ����+JFn���X�~�W\0����EQZN�20��j`#E�?h��o-�-��DSL�|�J����F,�	����;V�m!���b��}\��fp���ͺ�)�pd�ud�+�c�g/M�e�
�I�Ubo����M��}ۄ��\X(�(���X��g]��]~	����ͳ��KM�iΣ�o��Etު?g�x6��p���E��W�g+7:�;��><3���S!�t�~�p6#bFjj�M����
�Uе[�m��j�>~�حH��߱w�@�6S9}V�c��҇~P��8��e?�2_P��4�[2�y��aB��ƭ���m�D�7H�lJڹ�>}���6H�kƍ�\�X�t��оTފ��ă��6Nt��J���X��M��7I��$���E�T�+����k�%7������~Z�\\���>`�V�P� g�j}��X� ��Q9˒ ujW�y�;�W��B�*�@���`���_Ǯy��2}�h{bD '̵G{l�:Lsp�2EHo���{6Gk�]�d⓻�29�ႋ�{骏>tdg�F,d����:�wչI�z�ϋ��u
��u���uNQ#�SyB1V��!��c���8�j	Ų͍�[�2˒vrw0A�mq����{�^�ƃ��]��.7P:�`{Ȁ��/�my�|
d��߫Y�,l�-���2����!�V���'�.�L�2~���
==υ������ �L<놖�7�ێ�6�$tx����c*A8���!dݒy�)P��#��pI�RAc$�Ї	�Y������&��e�]����LT���<�C܉�R�9�ߘy���^F�'�G �#�ق\|Bm�9�:�ӟ�S7��Ҿ_`�TX�ǡ�~�gc�pE�s�
\Fi�P#�uA�$@y��W��JF`O|�~,�>�Z�����9����2c\��X�r�t�������; �UV	}���H�+�g����z-�����B��I���^1v��ؽ(�=���j&+v��9+�ܫ�[:���$��<�s>f�����?I�߁��vx��7Dk�.��7��}�uI�rל����`�nʛJŒ*_:� y��͂����`��ۼǇ�{z3���Iz�$�yX�ڀV2�sv�	:��=΄���(�M�Mm��B�R�kAb?q�ċ�����3<4#��5�!M�KI��N���.N�����H�	9A���0H�T1�=aX�����v�魼A�?�5�qwQ噤�II�W�x�P���e2�>����XA!2�yW6�/����s�d޽�BZD��*�i�H�S1�1/p�/�
��+����m��;!�V-���b�p�N��*׳���N������P��C�^���O�5��,�->�A���N�x�F�����] �|�τu��K�i��^X�:�e�Tl��,�z����"o/�y3�r�L���.%<r����r����&KM� ��n��S�M̶�ir.v��qmT[h�>�<	���QLi����i���EFYי�0m��ؒ�nJ�(�Z�*_��1 8�*	�&L�X�i[�W��бe�`�>{r���Mi��R�� �K
�*V3崜�1g1�B�{�5��1Z������Ug//��G? r�M�����yjʚܹ�0U�QT�&S�E|y�='���D���?�c��MZ�)��x���q���c�ǼL�;*�n��mn��${԰7�24�XYJ�?%�r�T��2	3�":,�����땒�E�@?��Γ��Qg'^�;V1��z���ݟx��q�T�ʐj�����|Z/��2� ����������P�"yHl2iJ�و�h�:����|�D�@����E���I0��cP�`��ڀ���]��`�q��ɒ�ڞFC�`΁�U��W����m.�ۡ���/iVv�~=i���S�F�03P�83�*�֩���,(�B񬻒�)��Kߍf
&����+z�Rf��fQ��޸���+��Z8����KV?��g˭�f��^ '��ʍ��u�jMѢUb��X�K"������l��:2Q-�StYBNꚺ���A���
J������bx(�����嵲B���9��馐�]�=�^���W���� ��X�%ɒ�U1���.�/�x��!��N��`���Y��E��|�_�Ы�Y���G ���+'A��ȳ+,�*Q{����a{J�ǚ�ux����a��vv+#
���?*q0x>F�i8Z�N=�\���r��`���E�k�+2����%Lt��W�̈́g]��L����.�?Ҋ�4��s�[����hl����[T �O�����1���w�����a�`�����Z��	��\� y���T�g��G~S��ض������/����6(V��w���.�E}�g#��n2�4� Ӆ\�5T�j���;�J�Uk��;9=�J��O%[����_�#d�6��[<'G�j�L����4��+P���z.�`y��"r�9�ED�j�Ɂ�f��Zӷ���=�����0���_\���M��|]�r��2� n�B-]z�U����������#�%�xr�ܘ��whd�OJW]Fy�}&�j�g���R����0{���Ot���9��2���6j�v�_�y��Eͫ��\0�s,�暦�8㳄<؞�]��^`M�2�{����6y��e�nH�]�������ݵ�w�yi�6w�F�@찕]���/w�����,b]��GG��'
�
�yՌFkv�~@� _��>�*���O�ʝьqެ�����^=��`��Wߚ*�v��w;L�l��.�2OA	�9��͈xl�#cc�I�۱�x��>"�<����9G��Vo��O���a5���ӃĴz"��u�ܕ��mDG�k��Q����30YJ����/�}q�5O�x�U�S�R�u�����.H��ѿP�Ԍ��hu�4쯞e��0�Pף�����L���q��h�M�޾4읏lȝ;u�ե��Ti���K�����۔�+?]��!}v�S�rNIXe}�eS{�_�������nwF���<��͋�������e���P�{i�D�{�e_�P�����c=q��;A��9p����z/A2�\����rz�Pc��mRc�|r�ax�Y�"l��w}��Ŧ�m����s��8���v.%�O�F�.��'���E�d���2�v�������K�rZ .�Z&}h9Mw&�������!颹 R
Z�¤�М��Z��(^ �C�/
�g�N���-���f�]Ÿ�uv�=��ec�������˿����Ț%kP��W/���юsT��n�ۀ���fP�����n��J�H�q�u��G~h$��:r� s�����~����3$�Łb-����A�����̿	���׈*w���M��װs;mZo�%j�Y�ԑ�:V�	��J
D�dO?-Y�����jiC"�3cw�|�6��O�/,CY�-X����?����h�������"Ra�����
��"m�%�^��߼q3Yږ�g_	���-�ue�^�TW��dӔ��������8&Id�bA��_�U·����h̃7��H�����=�2�����ꠡ#�uoh2�O��e��0�q	5N��՛آbڬ���9@�h*��}�(*�����O�g=��I)��&M��p��FZ㕉!,c� �X�q�(<��D�~�������nE�t!��fǭ�y�1��q/�,����]?~��bۘ'̿N�]�.����ej�r˰��|	EG�x�؅,=�M�,���\��){&�K��[�;I|.�4�W�H���I	��MM�q"
�8cv92��A�ߒ�v���|5{�'�o�ԩ��x�$��%%v�����!��g`66>�~ν��´�e�b��6�-)��X�1�)![�o���y�=$Ĩ��?���J�d���u^0�����7��)��9ɺ� 8��:/�
WW��r��p�{�MQ�����h�dL�t>�'�����
<P�}��$�ߤ[$�xՂ�E�M��� ��Y���I�.�-3K���Ei�`�-Dy<��RBvnmw�M��E�&���m�(c�z<�w]Uno������>�.뛢M�J�H�v��,��.K8��h컸8P��P1jRV��+��^Mc�˲'A�f2v'�sN��$Ф�?D!>�&�o)ǯ�脗�s\�a�������ܛ���(�|�~&�~�sl-f�=}~J��'������4�4��"��o�=���*�ƨ3��>)�*�f3�汌g��G"���`_i�t�[)��Ő2`�O	���e�A�������A�������Cƅ��s,*IW�x�,��YX���Z�e�새�s�2����@��VAW�e�b[U�A�%gkiI�>��7��:}���^Ún$�*�Ә��7~Pajj�<wh9�o��ɹ�����Qby<Ww}`��0/ҷC�z�;M����(9)�����W4+nXB�쫦ᳫ���#�+��.���➝&�y�A��'�k*������zپ�v{?�����U����jS��ݽ�/�W��7.�Lr�1�����w�G��e����_-
X$fda/�d6g�ͮ`������oy*��hp�u�v�;��n�L�%ʾL��zy��q	>�:�~O�����9�
g��/���a-o�������nb�2����su��"�`!uַ�'Iy2>6�-{"��P����^�N9<wLjh4�M��s�U�"�_��V:G*au�� �*�D\P<O�0cՌ�x_�dо⧭(U�b�w~[�s
���X%�z �齱��H���H�_ׅñ��M!t�yt�ꎽ4�3Bgw�eJ�I+E��,8�p!{�l{�{:���d����@�Nq�s��GG�����u��~�C�=�m�˲�!���L�ǐ>�;��B�NK��ٗ4]c�-$]��א5��,&���ˈ�O�����ޖ�}A[_����%�WW��1c�|��`��W��&T��[ҽ߻=�����}�J')s�<E������K�-�Ejj嚼�Jc�lw�J�߿�����u����&^����5���g�0w�GS�U�;�x��<\�2��
:�����Cc�����f�����Ph^�?c���=/Ӈ�E�A5dZ	<3we��]��t)�!5��r|�[�� 
�_t���.^Ä�V2����j�^+u����O���~Q��I�V�j�g�7|)�;<,���?jNr�b5�^���$����9���d��BU�o��ҋ��dC*<�z)�{�g��H�i ���֍[��
�H�1��U�]܈���l ��CP�6O�-M�[���]�����!�,�c�����A&]CX�vh��_mD�'�f3?�A!��"��T�nN?��V���N�K���He]ψR	������2����Pͨ�$�i	ı�Boy�Q��~`�pA��s�p&|Ȉ"�gHm�O����B٭
�����`ĘZ0 ��VGR��\��>��"�߳�H���g���{��=Lf��'�J���-�����<�@�����2�Ր��뙇}�n�Ή�=��̓�8՜C"�����
�	[	[�{>���"�w�-2���5l��J��|�Ps�g��@���*�֩ss����Ϙ���U��+8N}�{^U%Q�yq>H���xM�r��&��rB ��l���=��5���(N��72�o�3��ٙ�#R~�)w��
���������ζaQ���k�s�E�"��D��`�_��"��(�M����U.,���'� ̀b�������{y�6��i�'���aMz��d$}�FRWv��(U�s��2�	�2=�� O;k~N��.v/HG�Ũ�hN��5S�
�Y@t�AV7� ���lU�;�!�k������<-��E)�� �iƘ���y6�͟o�H���	�nQx�&�wҒ���Rɿ�ɇ]~Z�a%�Fd�k�
sO��<�������=.�kl�;yK=۠��L��}9'��X*�8�T[�:���Ǩv�'^5ə�:�P��D�ǈ�o˖����ʸ����zJz���kͩ�˴�}ח�n����`�>_KIpZ[��9#"��J�F��ee�txϬ���*}#B/�[��L�SjI������L��������-��;���f&$
<�L<����������@X��BR�Ա{��64+��w~B�c���ԓnla�]���1�-�`g�Q�D�)tsJ6R�x3�%f9<�&��6�'�V4���� P�J��>��'r_��)�K�^�w�V����Cܠ��*#�ޔ������A�٧���Ʋ�1�y.����<�3>��Ԉ@U�Ǫ^e�wcZt!�^)���̆s3�����(�|WT�L�~0��$�'�P��13',kTy3��͡UKqe��՜��X����}ʱMp�qsCe�R���s���7���.}6�$s����y�t���(�Ɛ��P*��N�����gF+��Mޛ��ۑ�d#�%����h���2%�4����I�2�>d	����7"�	trk$���ኧy�"�����*9�3��u��H`�6R�MG�c^���܁pE��+W��P1VV[�E�a���}�
��Am�&_Y$�5�2��iE[Nj� *D�/}Cބ�7Jc,N���<�����M2����>�R�Vm�C���]��~�0{\C��x�����s��bR��L�}�G]~�
Oe���jjH{y��x�^� U������N�}�<
n���p�����
e��{qG��\ǩ��3f��#D��"����72C@m��Q]� =^:>�)�L�d��"z9��@|I�b��Ǡ�rH�e�"w��!�l;ZT��[c�ڷ�<Gv�4m�@����DY���i�ЬtG��]���΀��џ#k�,��Bl�r�J@�eWg��G���I�Xq�-^����w��&�����w�P��e� �w�	/+�z߇}Z��J驫�-p���g��U<}�Ue�_s�='(4%F���=�4�����ӄ�3��s�,�3��n����7�B`�D$�n�%�\���L�(�1wV
�_@�~]�#2P7?���O�-�6|��ֿ������p�[�uUU�?]]9	@Y?[9a45guv�"X�/C-'<wT�B�Aa={j�IOs����Pןb EF��j.X����}�I�X�5.���\�GQ����R��v�x��8���Z`4-cQc�ճll��ڨu��x �
9W41'[<����f���U@I�`S�IQ&���Ԓ��&��=���]��|d"�T�Xm��W��Q^�p~�����E/�^�=����9;�����y���2�Z��;���)p0��Q�nK�g���yga�7�6~�ԫN�}-999pj��#r�����q�d��G����#�۷�}�� ��p���O��jLN-3�,b����9j��jz+�v��1oe&M�`�o�e�'��*�N�]O���[��p��%ٙ��3��^���	�R�zn����BH='��~�@���~��ĩ��'�����t��e���^��D�K=d�S��>���,�5�aH�M����NE��`_4�e��L�P�4�Ȗ��k��&G_��Nņ�oH��\�=�&�I���Eڄ}�ѷፃ����8d"�C����{��e�V�Rt��ON�xi{�D*��P7�
1���9�� 3���K�P��ܝ穰 �
Y-?���3x�Ѻ�����7�IT@=�O��;�;�A*�KxÙ�}\�js���9�r�[���L�3���G����2}��E��������?Ɣ���k|��%�-�O�ZU�bp�8���k�I�yq�� =�-�����k����t�rX���-�yJ�2��l�C!H� ʕ���6�Tt
[���=�S9�S��i��>���T����o�e,߇�ډfkqe�BD���3��@)K8T(=\�a�>���a���c=��u�̞�{�_��`���H�2��o�ϵ��dr!_h(�7\%����_��r6�EMW��F�'��9�';�Y_Њ��ٶ:f4�t�֠T_#���t+�f�{�������/5&����,B������j�Ơ2of��d�Bj�,�fn�7�n��1�\��{k�~B�NNŮ�([R�4�s�Kgo5,ԯ�}��-Ɓ��#4�/�7��E)�fvvz���
�T�A��;Uа�]�_���W��\��^Byyy�ؑ��Y��S$��q�������zF�����+ԕ��rP�X�j�k���`~��<�I��_��\��iK,e�����0LXa�]�[$�D��\��h����}ؾ�Ƹ0�)!w?��6�%u~���F��?����W,�����j1�\^�q<�vp�aJ�iAaN��ѪYUR����`�ʻ���5]��!�s4	6o��g�"P��AB�tN h��h�4�FQ���0�|0�3�p��ƣ�0{�~_������U�i��R}(�ޏ1�n9��&q�ı�����K]X�sR�C^��!1�WLb���A	����F��S�Y{0Qi{��Jg	:Z�U��oy��ԉ�ޑ(b�"�%��������>��k�4���l��#c�d��r�V���.���y+����]}�_h�n�KE'�A=H}���<l���%�S�y�ա�&�K�"�J7�kn��y�ȥPŌ�t���o��_6��h���Y S�3��@��`�0�U���Q,�E ���O���x��g�Sl��l""%ޯZ���4������CP��L_w���BZ�.�Z����<ꡟ��[#!�W3�Ս�u X�dx�����a�{��H3��N�PIm��,:�N�X� /�o�_�ξ��hw�Q_"X�-odz�ש���0 �ga�a��<�t�,�\J��Zo��񵪈��-�eNk�$����ZbB��f��K�����d��1�w��C�u��_@Ҩ�	���)T�lEc�d$g��%c���<�m	Wx��.�����O5���U7�|xb'��<��y���0ʤ��#E�z	��װ4���rS'��s�4�Wݧ"�\��D&z��#�V���E�$߇�%��ME}�A���x�� �Ș�vXa��7��p�?*�� �z��X7���e��r�8�[��Ed�Pqb	����I'y��+*�K�N}N�5HOn2�<��|��}��0����C�$&Y����,l(Q��y*f�Ն�P��̟v���WҖO�� R�}���.:�l�%�ܶP��������]4z�|UIEu��?����ΝHYh�C��P��O\&�;V')xv��%�f{��m���M�t�H���,Ȭ�J�%�o'X���#��ny<�%\f�ƌ��q` �[;ڐ^��b�7
������YV`�]�@1pl���޸��m�Zj�e�P���>u��ct��JR�ƣ30��>H��-�2w����h�k7Ϩ�r_,�}��@9��[Af4
�7�D��������7������E�t%EO�T��Ͻ[�a�8��dOGݥB��<��?�f�/�&$͒ݷB!f�����+~Z���*S���?yE�3����W-
ص(�1��Pz�����_ !x�����{[��p�]T������iV�-m#��]j�Ӌg7��T�y.�g���'��!y��E|��N���� ��jE���k��ę`Q����q�,��M��v3���w�_�]��C����}z�{��]�d(w�܃�݃����V�~�ﰈ��u^й�u��0$r�}���o���[:%�`u�~�������Y4�S�
b�m�����8kp����x�����^l�6��^{
\��=j�¯��L��/���rw�>fP��㒺����"xb����գS�آT�KV���=U�ˮ��U�5�3��T����(Ӓ^�t�ъ�(�ɲ���%�4�_?�mZ0�$������$�O5���U�]E�����eM�6����Y*x=T�b�ra\u�v���.K�������*`%M3URP�~��b��������&rW�V�����e8a��T�斷D+�I�/�2x��un���$��v�ZF�^��r]����2WTǲ�@����7��zq}���H�01�,�~EIII�r�j��&���ƲI���yF�Pi�~Ը�,�cy��GK.�fQ�[�n9���B��+�J��C�/�|P�خ�O �+3�ތ'��8��)C�,�� %���϶�54:��1!`��m7%�fZ��i^	}������oV�]A�9J�l�EbF���jp��$I�����G] 39���suc̿`�B_ƻ|�rKO�������0 �N��C�4b�k��3;;;;��q����՘��+�^y䵐>ʩ��XU)ݮ��_�� '�7���D�\���1 ��#�V~`)��iLJ0���m4�X3!�8K
��G�xF139���"�h� a�V��:�ڕ�m�*s�֚?�V��ݾ�?>2�@���I|�:*5|m�mT�����.Z<��k羄�<>���I��\�N&��au��(#ߊ�S��d��n�ܕ-������
��7��u�w���`<���F[i�|e�U�{��H���;|����N�x�=�&{��2�
�L����DUs�~�Pz(���=�K�_u�����o�t��I����CUF����J3�I�N@c���\]�y*ɦ*\��}d_�^��{ �-k��SkwG��C�^ޒVt�Ut�ؤ�6�*�sm���]hèW�Y�ӏZ�����`h�)�����׆g���Ӕ�4N�au�ȕ������p��ka�"ǔ��q��㖐mb��<i�78��:�E_F�Ph�Db~[?�;�N�U����ӧ#P�	�߿�џtL"*]�	�V٩�o"
�[;�m@�������"�� 5鼓���h��<l�Rt��<�}��UWP)@�7�m%x��ѕ���R0V������7¦�j!3�J��M�����G��=��@o�#�@�](�M'ݐ��tB|�Rp�Pts��q�{���r�r�xi�����@M���n�q;�۱z�}j6�����N�����o^������Z�3�M��˓[�Pް�X���*�2�q�y���511�L':�z���N�z�)�ژ��A�Lh̯�X����!חMK�!h�f2��'o�Ki���U78�wZ��!�9���x�
���I�R�O��S&#��a���5�Վ��n��^�Z���&��"�i���*��8�E�_qqqPs���`=��7V����/�� ���B��Ï���{�bf����6V!!eP��Y����jz#��Hy��p��V4���1�Sb���8Qʅon{D�ϯ�a�K��G�Uz���g���Ѐ_�i��J/w-��f2�6OT�:��Mh$����^/�5աzOQ��/t��9������Vw�q���S�D��2�7�P�����O���S*X�	�K��$罬U�h�F��u���L�a(E0o�ʦ�h��ŏ�ϼ_,���U6������Q�� ��Dn\�K�nha��]�H|M���2�tY{����!h����kY:�ae�q�'�B�����:]3�^�.���i�W@}5>��#��������[�E���㽾Y�v��9�~TQu��ZP@�|��Ʃ>�U��
o%����500�8�ĉ���[��V^-�)�*j9�X�)b99J{r�W 4��M����A���
���,G��xF#K�\?�l�^�'��EX����ʄwB}A�@�y1-=���D�,�Ím���w�Ըuf��^ ��0��ݟ���!l�6��Ч��H�x��n���,�L���_O�s-S�[(��At	�ƫ���X�&{j5l��J��t�TI���>=��j7�v`*���l�[0f�G.�%9�l-J��K�����>M�&��AM������?%EQ�`R��� f��4@��c��N��+�'퓯V�akEkK�J�����F��"v~�)� 
���n��㾻!��n-���5r/7��z ���6o�a���8��q�|�ҏ��`��P|o�y�7N��mJ�?{UÖ��^��e��|��#P����
k��#X���˕k��M� v5��S��(0�I�M�z��%i���S��D2�W������-�����Y���N��ʂ�(ɚhM���S���U��N�:rE��r�O�����ȾIy-Ol�LJ����s�Oc�\7�^s�_P��A�W5&OM��r�ܠ�T�z9���g�w��hV~�Ȧ
�9���r��)"�oX\�r
O$s�Ûۘ�NfF�%*QWG)JQm&�t�CoI���!Z)�f���6K}��Է�G&ZL�w}�8㓒 JI�ɓ@��n���/(�O�r1R�s5�76�|��n��x��]d�����G��A�k�P�S�������
c�� N��H�A�{�34��_Zoj%����N[�Ua4+5CD7O�d+��9
�� BO�r�����l����g��?�P��s��o�	g��y���j�M=}m�^)fLk�F��r�!�r4]2��u�[��և�y���j�L�}�����v�EL���l7� �
��ff�>��59�c]�P�Ivc�
b�l��/�Uf�x_J�T���l��J_���9��v�>v�gJ�v�L������$Ұ����"=��r�v�$l�����g"}X�؝��g����1�������K@�Խ�$��eM�gM���Z �&���I���B+��L\m3TC���y�z;8�P#��_�-��Th�Kզ��^
�GQ3A~,����:��9�jA��ż����}[��,a��e������O��M	�9!p���|7V�r����J.����r�����U��S�r��Y����x:�t�sfQ�b��#��h2�������H��54��o��*��4d�= }�u��
[��{NZ�_��(ȘZ����m�<[���׶џ�
�-.ag��;�Q�1��G�d-�1F��(�_�l��X�Qv�%���;h�����Fd��4+*0��B^*��mՏ�T���3T�ZP��R<uN�K ��,)}�iR�0�i����J��[�y���5�����;�/���	��_����ݝ��(<<}�}���F�+G�;�c����� u���|������y+��X���r9��Nh�j�g`8�MnCrpxd�D8��j ��=�XI���3�����^ܗ�ĕT�g�tm �pj\w�YL��!hȦ��[�{Iy����*��(g�|	.!?�z8��;��؉c��$��?�������A�//�I�v���rs����.O�$�l����4cw��2��8qjL?�2��L�ݹ�ǍLl����|�'��$���e"<[�Q��Z|-/+-�%�1�(��m�$�kY�k����OEh�ym��0�B���R����N=�뉶�.��uƅi���p�9'�?��}oM��>q�fR������~|�EG8�r�ߦ�cY��t����Ih�}&��jP]��2��^_.��j>��K��6�+8~���q�(��uEf�a`)5r�<��QW�Cڒ �cTqq�� �FS��/vޓ�m��p�z� ����P#Ҫ[7"��w?�Xx��u�JA���h�t�)#6�
H���3�K��u�R����a�m�����D�U��ՙ�p �7>8��\��tK{J/a��4���_E�dP��=4rZ�Zt�1}����q��>� �!��!O�?#�o��O�V���0�G��e��l�yÂ��f�^�m���RFފ��ips)usD:h�+��T?�L��T\ou��ON���l��h�� }x�P݊��a|[���Fܬ�ɼ���J��y�����y&Dʖ}�2aS(釀-��M)�����xJ���ֹM�H���?Gh�7�c��O��"-�G��e�����=<�t!�p|LT|]A��۽�C�j�o��,�A��D��ā�-���@��>�э�'�V�(��=��#���R��W��m�K�x�j���~��l_�
�N깺s�睠]�`��l��>͢KG�+�_��m����.Ĩ�����{����)=mj�a��OB&����`&�;f֝��� o�NQ3B�c�|���[ ���	�����pO8�x���=;�$u������N� k����4�m�n/G�,��e��Up��Y�T��S�[_L�~���Sj���6�$�z�P����Dl0ەw����V�� ���h��Q"A��LPj?�4��?�4�F���3��c<�#�ſȀf� Vە%�"(~���2���nd[^f�P_�&�u)�jxA�],)W%�đ�d~���nM���NN��WM�=}���0�Dr
#oiݻ��C�Wj�\)��?�������6I�&�k��d��D���Ԅ����j6c��}�����o���!j��/�.1:�{�'X��1�<��3jC���ݔ��uErN=��r�[�ˡ�����Ę�5*Q�k@������O���*GBd3y��˲�>�΄��q��cPe*�]���0�-Ķ�P��[^���t��{f����^���m߭�KJ�d�.�+e���h]p0�5�({꣈V�ʓx�r�X�"Ů���K����hn�ո�vi+�vL�X�.K����'�d)��:�ޫ0�������?9dS��ɮ�tdD�讄�d���SVG����EQ�l99Ƒ��BV��d�C���]o���{<�'�^�k<���N��2�g~ӯh�qiNx��R�g$��>��$��37�#XMuIa�M}�Y�^mB���Yy�~K�ːӔ��?� x��,Z���{�XjA3u��ro���{���F�T��(�<�m��}���i+?���:����n���k�v���B�����0���o�,��B��`�=-�;v��ș�e��m^���-�Њ߶�z���jAȟ1���c�OoN��� �i�q3_e�0q��L���ֲ:��%���������},@�z���%|�gpp�kx8k�+A�4Aڠ1Y'Nݼ�����=%<'*T(44t�m��Z�s�q&��	v�ƺ��p7JN��9 k�Ue%{(��� �t�Q=R�6������q�F���� ەo�ׯ��jjj�_}&�8��օ͗A���33-w9��'vT�~5U�q+mK�':��G;h��J��=��m��)^++ny^��M�����KZO0��s-n�ЃNyq�"K���_g��F
VPWW��q� ��03Lޓ��u�EԚ�u.W�Z
j��OS�Z�0�jLLX=nk}=8��u����2��������wɑ'^�|��e����=�%txE'�<�%�5���S5�����Ur���nCӱ�A~▽VXQ5q�0��sm'"x��˃�z�+����H��X�nl<���}a�޳ۥ��y��l|Rj��Kv���k�ќ�S��a~N��-}��:\37�X�#�)?=n�ٮ��p�F��+}�J��7&�i�􅋕Y�Ž�ѐzd�z%� 6��U��Ǧ��iȧ?�7���I���Sտ�C�9jUA˼{��j�%�Ec`_?u����@�7��"�h�!����'� ��$rL����#ZI�^����JW�N�a��4>8��W��A��'i���NL0ϖ����b�j97�e�b�L�����|о���(]"��S���p~��ku�]%%Ogg��С��̱�Dm��Pm7���{��W<�OM1��Jc^��$���ʲ�'��g����s�R�!����!�&�G��j^I��O���b*��ia��ӳ�f�%v_Yʟ��Y�Y�q��u��ͼ�b��]O�ۭ.s�6�555��v�h��\/��EEY
�m�`}G��'Y����72��yE��8m����=&��x� o.pM����P��ɦ��Bp:o���(]����w?@II��zr�I��tD���/)��+�}���}*�49Z���]���(��w������lV�`�A#%ޯx�����UE��N����Ӑv�=c��J���H��+�����D�Qć�⯛����C�I���J�x�z���>�V=X�#cxK��XS�
��3��RN��`���NE�U>�F�9�l�)֎%���Byu��*PVl��ȕϚ�z�h�c������'%����	�F�`?3���e�p�c���5�ϲ�z�x��2Tߨ(�>��������+?���k��S�E?Qǈ�V81���!9��z��v����z����ыd�2)j넄��L�g��h��
5��i"�o*d]b�N�!G�Dd_��x�	Ý�;����$m׭�	{�VZ^~�2F�� �|`&�yM�N�Q.4�^%_�F�7x�x\��/}��_Y��W��b.�[n��R���]��(��瘖�h�~/�w��g�=Ŏ����?��������,��OM��H���f�)���m�Ճ�|���Cᒔ�]�����6=+.Zb�G:�F��_#��. �C����x�f��9i��9]H1	��?�������1��=�> �PȞ�*IЗ	\H��{�cm+I���	)��'骺��UUn>�~qXwyk������������Fp�]�	i�r�Y��-�Я��x͟�������t�dW��qT�� �ɷ[�J+** ��~TĒ��K��7��D��Ԡ`kk�ãzb���`SsklD�[�34n��l���O���O=��l>��q����g+mi�d�jƏ
�>��u#�~���'�˴���@�ͪRc�=Z���������_�ml��,wz�E�`'C�&o�A��p3�f!�h����?`4^����'���iR�Q$ԭ����&v�+^ԫI�颉�Q�0r����>炶�	y����a��΃lD�)� �2�&�o1��2Ÿc�ֿښ}��(Q ,3��ۛi-�# G���)����Q�V���M��Y��Rl��v�==�Ū�K�A{=���0�*-t:���,U\.�H���a߉�J���"&/�Y�u8ꘙ`2%�?;��F۵�X(�,��t���QV\L�� ��W3h;��í��W��`�w�$�u����@Z^~S��9Y6��Ca������+L���f_�L�W�c{V���ܳ��&��

�֏����&�ߓ�X�������'�/����T�ѻ�G��f[��.'�/6 a����M���i��Vud�}a�;��&ݣ��зdt��|3��	�am,�%�P�=4����vS�o���ʰ��j���85a�@_��֦�&��m�ǩ����X��[iVb^�Q��
���hN@r\i��d�5�_�S������C3�����i}]+56�B��z/�k�]фl����OV�:��\5a���ړ��l��0��0�B�0�_JyM�@�qz%=�JF����vpx1��E��s�F�qvmD&P(7$��R�	h==K��~S�Ԫ�m�f� ���J�9,�����_���S���vW�R��׫5�$e�t���񲲱au2���?X���$�<_����h7^O96�42RN�iS� �D��3D�K#n�f��0�[����ֱ����wA����y��>�'����#0��$�������r<q*�>�2�GX�M�/n�>0O=-gQ�}�ڵk���Wն	@�$��Ss��2^��f�[bp�*5�F6vr.���e��<�u�H֒	���f����e��Q����TK�09�<7�^x���ԯ�ȫ���	�_����6~�Hz+���A`;6":�7��8��e�����YZ���[֨y�r�~��o/a��U(�O�y��7�ۏr#oHE��Q��6喅97A���k�N�@<��i���8b�_�����F���>" S�K�G����/��<�8s�!$�Ԉ��#2�~���;��ȾT(��i���+�#�0�T�2;q+`�����ܜh��r|��4�?؀%b��$tv�$&�͘���uԛ���ܸ}�v��[b��|&,
���Q�|��sk�7����2�?�йq����ʕ��6"a8fO���E��.���F(6���j(;�f�$n���aᎵ]yU�b�L}�-��,�Аkn����"��+�.��*��u���3�U��?�ؚ�32p�[��r���b>��R&�<Y�P��G��[�O#r��J7�^�3�pJ�/Mоw��%EE�����͟{~�2͟���6X�+��)��nl�Xm��E����j��K�h�dLFj%j�4��������13ށ�`��`����"%����҇;&�Px�_��V�?x-����W�� =rn����NQ�A�}	���aGBr97ʁئ�A_Y��iKȐTza����Ċ{�l k�*nO)�����a8nLHz��-�]^�vw�F�tPj�r��۰I> Zzꑍ����!lp�V9��*�؍� ) ��z頋�N=>�U�8]t�od�sq`�ݲ��7u�����;_k^	l�,��˃�tuoFV; q@��p7Z�����l>��>���0^�U1 }v�W[�s"Ƿo����w�`�����f���l��ӣ��1��	nA;V�nx�R5x7�������ܬ2ʽ �5�Ǽj��dۻ�a+�U/�C���Wf�Kʦ��I��N�e�=Ы�֏�.��>'}�Nl�A q����θ��&�B�w_�	W�"ޡ,&���|� �bs���gI�߸0P��R���&V&�c__@Ӡ�+9p���0��+�?N��S�������2C�ih�ӑ#l�7�n����c@������� 2��v1��Er�S"��%�
h"3��5��y纴��L(�O�ssHC�w���2�?�;dWZ��ðy�d`���%4D/��#�3(�)�%��M(]@U��]/����X�xAB[�kVV?�5�Q���b����
�
ac���4��I��Nzaha暎A��IX˱��}b�6�z��qn�0��<7��4.��H��0�}D=��R��7�
�^ �U,�=�m�m���������K���OT�Q[�k{�5�qP^Y���-u�[.�F������[in��Y6q�zdfhtD�����SH�_g�7�,�gJI�/^�|5&�`�����Lk{���_�0�2i��eI�vl���tU�GIc~�`O�Y�����p6@E�C�����C�S�]p����(`v�H���jLM���N�iY":��s���3a��i��_=�*�7\\��Ҷ���,��#������I�9Ɩw��l�VSgN���?�z�87D9�#]#�g3�e�+��B5���^l����n�_��X��f&���ي�o"N�e��0�����8$��}��y�Y�d��=,��e���vb̍�0�S^K`eR�\�~o���F��9�g�B�#�pz��<񔀂"P���~j19-�P74�n$�^�\�s�����--iZV�AbY-�4~3b7.z(s���ׁ:���+�R3`'X�ĚFG_������/;��4��ɖV��Y�6��ne�V%8��C���[W��ސ�X��T�&gg�� M��TVT|ו#P�"�N�ƕs>�%��Y L+)YH-���T�i��X�\��ȥqeA.b��n��E&nE�1�K�[�Xoؤy�X��jKQx1��NSS+(��ƹ��v��S}��n����RPRB/��J���t^��x�����Ye��Ҕ=}�^��ުl�(��NVfwK���@�z$.T(Џ�a���>(���uh1'�2_tm��P?������/<3��}�Fh@}ϕ�������Ձ=��:;��OҊ���I�
3g�1UW����8K�89����]���L\����|Lo}8(&�}c Ia��*.����n��u�R����vjMxhh:�QA�u�����{�P!&��5�vևրQ=|������xs �� 5��k�}O����Tu����S����ӫ��t	� w�t�t�[5��{3�ޚjSc�P��E�2��΍)��f�Wi�!�ӏS�l�cx����_�ul��O����?[ݍڞ�db���T�G�G���Ɪ��w��vWߍ��H�s{e�s�$drf�z`��u^I���j�;��bb���������7��45e�Z;#(���K�f�����{�c��#�/��ޮ�P���%��ƲR���V�(�����y3֜��s��H�Ϯ�n�d�92�_�~��s�'Q��G�[g��ԋio��{j����˳��:1�̙�-��d�v)���f�-�WJ
����:iђ`����tǽ�ິ�Sd��U�����2H��M���1P��Ir�SiZ���r��r���ai��#�j{%���Q�t���Co�H<}Z��6<��vW���,*�>x��2!�������C�+���;�m�˹���6�B�߮q�m�j^+'�g[����/�z��@N,M3�QO�Ac��>/"4�p\��p���"���~0�c�W��cg~�LVĆn��\�^��Z��9���ڍ�g�Oas|
����Yp<�A�9>Å�&�{�c�gN��h�~p3�����+=�a���̓;����a4����z�7Htwt!{����{�]n��F������kc��Z��c^ ��\ �1lm��C��\�	��k�=��`i��~*�T��5�Lpx�F��V��5J�p��\��\8��=8�}DP��(XN"}�:��6������Lq�e���r)Z�z�}�=u!΁���J�|~��ծ�����F_d���w�P�2kl@�v�YE�N�E�Lp:�ʸ��6�x�?5׻]���U�+�~[��&�X|�i��JoyL�p����{�O\�(��XD����1���?��uߘ���.���%���KHye��}]��xYi�(����NǶ�R/�nd�|@3� 3�z�M����J�Z��9���H�0- )��S��4���O+9P<Ի��À:gA�O>v�����������L6+~j������'w!�c��W��C�7������\�N��0ڍl"�#O�f�CY����a���d����~T�q�vy^]�m*����Nݵ�"�jS�T�LM�lO�SeUϬ�/>M��ٺ�.��׵�m�������u�YW`���!��f�BBDGL��0�^���)'���k
��<!ٞ����D|E���u�&�|�%f)h#���[=��,���!%�e�`�{�Km��0��u�3g1�25f�1>���h�ދɛ��y�Wd���%ج;6�q/�:y�	�N������֝�(�c��{Fx]��x��N�lI�<���,�YZX!��n޻����U���cS��M������{*P����N	����v���(�a�W?t��9�Q��,���W�������9�GZ�m�KD�M���!�t�lRg�݆��<%Eˊ禧
��wK��/T�v��i���z�*�n/u�,�����;�Ζ���>�hi2B�_
�J�[���Қ���?\)�s�,�u��![>t�ݘ�.�1P�E7��Q���A4�לk��7B���<H�%w���A�-Iy��H L.��:�\�M,�l��)b�;nm�jH�wePÎb �Z�Y��@����ҳkՍ��������:o�]�M��e.��Y��	�B��5
7���'�m$9?��~]^&<?ϢQQ�J����Klu��8ۭ�xD�.A?�c�{�@��WF$7���m��Ŀ=��g�������rU0fĔ׵��*����8r����yv�gU���u�'����V	�a��\.�do�����<�V�|!$&�U&\��qA�W�^���忱x���!�����΋��a_U������v�'�\<1sJ}8|-'��Q��ߐ�2�))lA����v�_'E#kj�SQ�/�Gb?�x�4s�w�
R�eqrph�%��s�j��g�_Oˡ��+����7�x���Q����#���URY����C����{��ث1�X�-! :�n���SU�V����u^�Q�,LCj��M6�G[B�j������ݏ��h�x4������n��R.]�q4f��׍��3�,���fM7%rX�J��s%&�;��]��H��+)a�]�a�Ar��ʏd�zZ�f0;LEM���=�c����� +�Ia[��d�O�����<�4�&r�ˆ��x��Z{���$W��
��Vv��B��ͻ/9c�ٻ�����#�'i�8ɫ~�����JOǙj��E�'�����řN��N�`�>��ؑJ�b:�[��;0�Uֆ�84S!T��u�XVTR����k},*p+��S��s����n��Q[q��\+'Rj��@���>����g,�J�%�
�Ŝ35�t=M���,�e"M@Z��;�+hik$�l����l|։{|�}��`�o�joK�Ӯ>�wX9K����QN�$B���ѓ�a������[A?��b���2)���:�C^�%��	ti��W)�m4�J111^��GX￧J�Ȳv��>�T��AWW� 6J655a���|������z�nd�M?�R\�	�����?t�N��Y,..�y�pa�
�����5'�����3��� >o�)uzĞ����E��~���;�βݗ��Č܋�q��LfG*�>�	�����w������&-��%�,��P�?p����ń�W��K몧"Y��g{y��Ps8쐙KLa�7CCM�@ch�+�o��-lSB�u��F��m���w��YEf��K����I��?��\��k��_���۞&���/��������;n]��D��Ǽ��3��ǂ%�<��&@W@�U۱v�kR� 뎮�������#�H�� ��aq�Px��X,��' ��͏fCa���G��B�3��~�e��&�����.�w�p�W�a�XE��}'B��'�p΅��F�W<�ǣ��u�	��Ӵ,E�T�IK�|隋��չo6����GHK�r4�P_Nq��RMC��~`���}�����sU���fl�:��7���ފ#�+��N�
tH���C��|�B�GOlWW�ng�
> ����Ü���>�j��#�HDw)��k�FK���1�|å_1����iPc$%r��Ng��+�r�<��F">Kv&�E�$BS���jv<���N�	`A��-�kE�Va��b�[2�u��Qx��/�ѩmv����I?]���ƤB�,b/�\�bJ<r^Q�(������.��Gi����4������t�0�2]ӵ[�����6��n��������s��?3��!-�i�G�Q�3�D�۬|�7����0���Mi�[�Iy<�,�S$�O�F���	�9���LWV�d�-��[ ��GOZ`��w�4)�y�\7EHk%m�2;�=�ug}RZs䯳}+�程�
��C�7H�jl�J����X�'�Ѻ4'�LN�(�ܯC��/,77~��E#5D�~2����.�b��!�t�f��F	TUlJ�*��Sb�ώ���f�m�i�A�КNX�U�9���'�Ze�}�/e�BM�u�[�d�dj.wG�MԾ2��>/V�J8�K�������CZ�^[��*\$�#���3�ϩ\j��_)N���ש������WYe�8����k��Z�����NZ��V�������	I��6��v�L�]�C�v���S#��7���8�`x{[�;n� ��>�� 73c⦟�g'��Θ����X���S uY:\�&���iݫ����J���!��[���S����џ�_�u�����Ɗ��`Z���D8��	���1�[���ڽ�ne��0ioY(����.+�t��Sct��[���}ԅ�V��qa�X��{Vw��oUX�8�bX|�r�e.����y���n?M8|������V[��=�d,�ޯ+@��?1�,�s4M�A/��9s�4#���WEA!ܾU�A�r|����:����/�	{dʽ	�8���:��)�*�*��g�SS$�{@�c2=h���h�|���VR�B�0?���ز���wa����7>��<�.�6';"����a�\�m�n���OL:b6�0���lJ���5�����ޞqįD��6K�/l&D��)����:��0��~G�4���|t��m�w�g�.�B�;h�  96M�S4���cy�1��L���a��GG��CI8t�����FM�r:@9����wV�p����'�لL3�B��lӂ�5��I�Y^|���� �Č)�f�u�ߟ�̬�;���%+���)����9}�wy����0�`�9�9��F:�K5��zIfKb<Xq��H�٘���Y���q$�m�+�e�?9�Z̟�9�PB;k&��r<�CĆ��Ѝ��[�&�2��.�Z���;��`;�sO���7]~ͬ=�[X9Zמ9޺�(���)(`b�ګ�~�KryUPקE��!���1��I	��I����d�#�v�H�ॴ���"\��q�� *~=xS�:tb>�ku7�M���D�u��?c��[������>��A�1mZ�X~�-��5�Wt��8Q0�����ҷ��'�����?�H$)5_k�on(3��:�Ǩ�!��b�jo�-�3��u|~vl���mf��X�6���o�f��d��S�Ҟ9������l�Gi��oi� ����an�+j@Q���iH��zV]~�EN��B�Oݺ����cz�H�@��I�O,,K+x�{��"��ne	�����6�*8�+^ـ�S+9��$�ZgA�3�����J�.VR�v��9�.�R_R���R�A�uj��D��>F�TW7?���q%��o8e�1��}�G}e%:� <B���y�L`n������~�Q$�Uۇ�w�P@�Ը:ܩ�����(����J����aFc�!9Po[S�p���Bܖ�4ŕ{�1!/�+L�����Ջ�:q���V�T��&��&��g��U���ׄ����������g�u#S��*�@7)[�݀�~f�ObE��(��h��y;}4П��+��o�3s)6GA��������̄)�6�o�5ٞMVJ�\���(��)C-�:�U0T�����C��ּ{I⽫�_��4�jeE4�]��լT����?Q��	�����,�A,��K��v��1�$w�mEb��I,N'������ �K�"�{n�(7)�6�˃�z�LW�� ���&�_�đI)�o�M^?���O�%y���G���7���H׻)y�EIl�^���DM$Em�"��F��-2�n.��C{��&
>�~�b+od�*n-����;"H}���ov����g�Y�o&�y6�����q^��]F�U���w����V�1-A]�����S�+��y�xQ$�o@P jȼ����Q%���u�s�?]K?�t���Wc���w��[en7+��I�_�����R�V^!�쥙~/��4��&�t�:��j����IT��FEEř�t�}��QԷ�R���"{A�j=���-.IJ������1�Xh���Ť�E�1��ts8��5B`Y��g��k�x��6����y�����a��ȿPUP~G���n, ����y�� �"���8����qY��4]��P�����1�P6+��;��wZ+�O0�����"�z������;�F	���Z~E��!4�2�� ���*���T���FB%{a���ȣ���=DE�V��K�W_�k��_�mhOt�n���Uٴ���:��%��q%����@A�UnУ�
J�LX��K(�p# ���S�b�����Yϓ,���f�R��֊�W�n��:�/ũ�dBW~����	��Xz����.C���g��=p�(1Ff�f^�ҷо�/3k�AB�md ��2�E�Qи:�1��)��f����P�����\B=<�t��D�y�m��D�ʐMh���~�]�"�#���X�_�ޙ�E��N�ܮ��8��K�,.�`�%y)�25��|��e2GM�H�mB�c�=���Ր��(�f?M�<�s=���\���aQ�[����4�����Tf2&��<f)�7U���bl��4Ѝ�����f%�s㦦AȺ�P��_�M��d�߻����fe�C �y�y�%3�阇E�ܹ��;^ vOW�n�ΝD�MŠ�y��ʈ���� ���;fD=ۺ��W�OL����6x��X����ĝ�]�=���s��R�9K�/t���B�����:5|��:,_'=���Wt�ǭo;m�CN*~�	��3��F��T<�$�gӦ�Zs�ܫƙ�r٭4������t�F�jc�#Il?�t��@�2	�O��������\8ﴮ��焯��Z |��B�$-���1*�hE�A��W#8t3��3*�BV��9�ʰ���R?W���u�I����.~�3E/t�z��m�sj����!��Ԩyq�;h�'z�� *���a�����!��~Խ�67p؋�K��������.g�{�i���;�_ɱl�
^�e�ZS�4}%���dO=2� ��~LV���V~����5
�*V��4����=�&Dl�Ww8� <Q��$NͯP]���n�>��+`�>Jz�0/;�c�Fi�=ˉ�|�:hS�k8�R퓝jU0��l�J7��j���{�x�z��� 4ݜ�z���J9�s���*�����~�.V��������!)��A�1�O)t����Y���E���L�g4c��`�g�!��Ѣ��gZ�+-��6�d2�ئP&�W���ș�R̬R�@�r7؆9eĺ�	�M&����8 t�nj�
�0K	~ڦS�ș�ӧV�� �֟�ӾMIk��}���Y(�^��G�����Kn�X6~U �o�`�V�0�R�P;�k�A�<"h-��ͫm"ٴnJ���J\/����"T"�^�&���SV���M�z��Ȳ�&љJ&�Ն� g��B80���׶Wt1�G�g�^іm�AH����ٖ�u,T`�:7J�̖8&P�K�6~��*�;{c��NP`YSǯ*}�es�	Š��Y�cA�$����9��=*��J�����O`����~Z?=�j	�-έ���F���� +�J����mm�Y��
z�gP�8��KD�p����K�di :��)�_@�3��t���g��G��_K�S��R�]S��{<��&K9��ݐE��N����4p;��xb�21��Rڐ�6�W�U���ՠ��#�3R��0\���G��-q�B�1�[&�����*İ8 ��6(�|�a������1� �N,Z��ǹ�Z�-�S��=! _�w��q���V%��O�9�
��}�p�u������&��yqhP'�N�|c'f�4�D��������#G'�_k��D��cP���; ��ԑ��0�ʕ����rm/�Y(��oefV@=�zC�.p:To�Sf'�$��{�T�P橺���V�6�D�����xF�����H �Ǚ�4j@���ȫ�l0�����PasLI\
�`eflv����<k����_
r�0�艀44�˄k�>.Ëߟ�?��dҝ� %�j�i	���NZ����w��u��/w*��a�����g�݃��>��������/�0K�~�Y�Qk�^:�n�_\3G���XS ?�$Ǘ�2�Җ����ʹ��DGr�������?r�ey-:w��Ma���q�[�_[���ɑ�^~W�,�ѻH�1;�}`@s�m���p�� �-m�t(��\?��;�에�7���Q���f>�	\w.��t}��J�=-�E�L�����a _�:��������c ��u�����$'�N[t���<���E���Ō���=��ro7F�,0Q}�|���A�������~��v�w�a'bC�g�G���cxi	�y��s� �8�w�� b�	�?6}Jz�*H������T���lD��=@�PF6�ȩ	lQ��C�K�j��-����p;�u���H�b�gL�&(=��G�����0��D�: ��q�@�����=��#��GI�8�_q�Ys.�7���RE��h���:���_¡�q�SS�3�;п��}�Z:7`3�����(cr�[�@�f��/�����v��G�s}�����h����r`�(&Q��ɱ�a��0�@ >~����Y[k�]��%��.��%���',�-��/������A\�'�_����A�bͯ��J	J��<}_x�ȸ؉11T�i	6��dӼ
+����
|/*��{���/�aϷ�tT�s��%uQ��CKe`��W�G��|~�}��L���=�ؕ�N����׻o�|@�@���J�i޷�v9�7�ԅ@O�tr;
T�>|N�LE|�x���_��C�,�v��M�gdPHR�&�r	��.�{��ز����y�N�+=�N��8���_�S�ܰIwݿ o]�N�+cb�_�3v�Kڧ~�/�1{�`��Y�Nr���.ՇE�eڱЍ"��a}7���B����LX����.RP+_H�f�������N��2 �.�3��a�Q^ϛ�ĩ;���㥷���O�lTr
���rf�y�:I�ΘcȄK�
�S~�����> ;@m�	(��bJQo����w:�S��U�f"7����M���=��nS�X{�Ӆ��>�"��/��<��Z�;�q�����(�wcP�,���Q�An���I�*�l �P	����J0��=|�$��d�h���ǾZs��UA$}�ц��-y�p��(U�;/z�!��@��G�ʵ��2���r!��p����;����;�*&�Lu��2���U_�z�7��A�v-��L؛�6׀~}�*�3��AJ��,Ԋ�s*��c�AuN�f�����۸P՚
jc�j�3/�ʄ���I)�`�u�t�����"f/���2�D���8 N�������j`�r���Z�t���F��g�Kb�m fRϵiJ�!̎���~�p�7|-�M��b��L.�Fj���^�6uI��Zf�[�ָX���@�^Z���<}�U�Z�˪M�@#)8݆�8k���,��Y�|GNO1V`�]M�2�Db�ૺ`}�>hx��>k�Ʊt�-IC�Gq�N�$Г�Tgi'��a���� c�I/T���/���x��6��� �٩����m�BR�>�(3	��5���$�^6���w��D�ۑ'�0�����
�pERPyL�(�D�65���/C�$�j�
0���J)����߂�E־}y�R�,�KJiٿN�d�g���y��s�-!�����^}���r��`�[�1�e/���-��7VX��0v�{u9o��?z�?���8ٵYa�ͨf���p����ӆ�l~�(gmI�<��>��;
��+P�i���a44�,���U����Z�62Pu<1�|�i��-�;�/��R�@w���4�w��9^9�M���B�2�s��
�e 7Q��Q�U)w��� pF�`�����]�Z����� &4�ŗi�l��+K�F~�{y��C�-v��y̅iMx_�k+��BF�u�<�q�w.��o�=�@�U��갾Q�W�Q�8�2��7�g}���$�.R����U�����@$O��Z=mt^u�V��/o���+x�l"լ�wI3_�[�Wԣ�/���+_5}�D��C�$����▿��Of�(�u`#n�O��9��W���g4�)��2N���{*������X�J:�����(�d;�J����'^;z�K�1�~�� �Č��	��r2�' 4�c�$q(����#�^n���%�Bhjن�>�ϸW#��"i��c��������5J�kJ�5�(y�6-�f݃�W�cb���&��G��J�m�Gu�)����V߻:�=���v�%��#��6�KhK	� �C�u��85��u���{	_���ɨ���H�^�&]W�/�-=ŧҤ[l�f�:�i�N-f��GA~q�u����7�]i��I�*�K��M~q�^#5�t�������	�y5z �@� ���t)(�c�ێ���j�J�P�����oB[d#8LׯH�⻼�8{�I���yl��2˒��%E&�o�oK��t��ޮ~X�_z�8�|�d�6�Í��PW��1\��h�۵�漦���\�)����w�_�c�"���B�va:�� �2�W���';	�~͟����
5RE�dJ�����ZK+��`41EC�%ߺ��k_���^��1�D����!�G5�͑'`hs炠3�y�+l8۱��������[�/[v<�!k��Y���T9K�k���'Ǆ�x��J�d�8I$�NU�QA؇Jd��6�:6�����(�l���}��n�W�l�JVOݫS�n�Q8L�K�&ĔA{����|A��
�>k6�VLNq���*����x�#���b@9���*����i2������<}�mF�ة����U�'I��#+{�L�P4}�+�������268�)3��:(�-!U��^]RcC1�F��lƒu�$��N��A]�������D���W������S���BMw�/1��I�I�'h$�|:鏁�����G�[������@�O��~δ �Ҫ!g� �4�Q���~F��/��E�\�'�W�),���J�2�u|�Q�j<�����͜9:L7�)U��	����5��/��}�ⰾN���UL,u#�'n�g��g�[x�o�ˇg�m:�OPq��Ԗj�DY�����ӡ���� :�����q��
�r���0���[NP`�������"~J.w���)>�~�XpHeZI%Q>�F�%����~N��f�hx��S	��a��[��|0ܦ��0�|���c�1*B�?�XJS��,�/FJ��Q.bp��$�8=���h��i�oD�σ�$U�.  �W���b�� ��FZ��O�9�=
�sʸt{A�'	fy����O�����a;�&bX�{�-��~�#({e8̃J�!�r�P6;�@���aiQƜ�FxT�����v �dw N�}a�3�6���^����
���%���tM�8�6��b$  �I�V�9 �F%X@��E3�%������]�DY��J+T������S��_Q��1l]L�e���;�
Eנ���kDFj��d�/Ϡ��@��Ρ!!�n>_���	�r��5]�H��\�b�|�̢(�0X�S�s���F$�`2����{Jk�ʁ[6��V�zH�y�=��QP�!
� ɻ*��gb�-����-}�?�DGX�oc��
��F��P�W�o�h7�m	�e,�b�k��Ą�h<%�������ʶ�<Q`���Z"/�Տg�0^�{���a�s%���l�������Q�P�"�ߛ�R�
�լm��"y9A=�@xb��
�;ٶ��#�y��,?�r���lBS��f��9J;��.�k�埰_�yf��\��4�g=s%���
,�D�ԻJ���d��m�1N��k����k������;��~"��6��l��iD�}!�qE�����S��5�����V���ب�A��%���e񺯊�YK>��N����D�����B��(�14X���Y�i6����F��s%{.3ᚏ��������0�f�+0�~���:�9����D��\�#�R�?w,�j��l�P�/l����|� cA'ЦG�{U��X�Z!&=�^���\�,�WH�Ls;9��w�Dn��sC\��LH���Bw��T��5��H�4�J���r�+x*ܬ#dl�,�S�k!���_a��O��5�S�"}���vL�	r��ï�R�������P�ǳ���"�E�{��i0�A��=��`����U�59KT+�H� ��0Uf.��#3	�����]��F���P8���/��{����%���fC�ei�}ɾ�]c�¨�-%*#�d#!	E�6#K��}_~����^��ԕ�>���k��y�i,l�E��p�h�:�Qe5��4�Ԋ?ߞ�mw*�t����mM���DYfg_���d����O�u.�J���'r������bA�A�js���� �Ӏh5�SC+���ʟ���8���Φƫi>H�@1ʽ"Q|����k,,�`�$�� *�ߒ]i�ʿ�~J���S�м3 �YF�+'�����`RE����>���H�f��B� p�;��Bo�vwQ��K-x���92w6�Q �,P��u���K��A����i�)!��C�3!�:��+��nԠ���n��ݷ�?9�-!��;43m�s�V�.V�AJ�;�"����]������'��� ���n�*��#�S�M�@��Op�Kp@�ټg���nnZ�w���/���3xV,x�fyl�-��R�����L�$P.�*s;�{s�(�s_@o�b�����&\����}ޠj	{Z׿�ê�.`��w7��{l.��ć�,C��O��c"}80�aնH�@_���xm�A���|o;$Q���r�R����'�
��N���sq8I~p�P6I��,@D����7;)�^���r��u��y��Yz����Yi�awO=D�P0}\/G稙AV��VS[����n��J���]�*KMBI��9��LJ8]���<��31��CN��N<
�+@���Dۄ�|��+��m��7+���W$s��W�5WQ^�ʹ���A��7\���Hh���f�d��^V�qm��^~ {}����T�+jmQ�<��'����� W;^�	Oɾ�u���jw�m���1�p�!�+��#���Ns��'��;z�s���������%���K'��{zz S��P�K���"�7�i��q�ҽn�8%�7A:��M�j��!�:�;��*��e!SU�	\��o�9f���)���u�c��R�#3�oF� �8������@G���-�ꑀ(M.f����3$UB%!Y�C��|Dn�	f��j˭���왯�6��a��7L�DlAy^ڿr%�\.����|?���Jc��M<%^�m�^�ؼ
 �4)�a݂�FN}N����a��f�9h+=�ҕ�(��R��|>�*S����ࣰ�\�O�{W� j!� D��������]���SBJ���,?G�܄���'�ɒ�ơ+��ӫ�n2��������"獀�����ujN��>�ۍ�X�4�.To�м��r&�M��їV��*tQ���@�e$k�2��Ea�j
P�q��y_����X�{-f0��c�����x	��ᖼ�eEM�BJg��!���֗i�� �~�$�R;���=����'?���
�>�����|�j�Z��.Q�D��R}Z�͖'?��>�,e��&
�+˛v���)n]�]-�����D$'z���y?<_x��C�X��]HyEj�2�,�`6�7��mM�����d��
�e�4���ܦG�o
�=x��r�	��TN������#��@=�r]L�>/���X��隇���,�QdzUϸ��e��@ ���������u!��h]�0���"��	J�zru�^:)J����|�f4�g���ɺ��W��,`�⽻Pc��NA=1��ح�����'g�O�@r�T��?���F�?�~�@�b�=�T�6DKL~�Y������5��� �F�ų'�e���ϟ!F�=�T���P�:���{"��|̃i>j�Rb��m�}Qjʗͫ�P �
�J ��v0��2r���;��r[bZ�@�e��ua�.�ToQ���D�l�Őc0t����jPҋ���&�d���!�H9he/��`f�s��>�8�/�,��?m�FhO��D	��v�����dʔyv�/�X��La��k���_K$�RV��x�IYEW_u���.[Z���Q�3^R�$��]=�=�҃`?���̾��3G���P�;/��f�(fiN�?SW�%N �j�����^�d_�5F�1�Rs G���S����9>����,���y<S�QKՋ��yM�FMsy�;'��#]3�7;{�u]�:��3_H��'%�k�\�t9�����RF {Ӹ#P. �xx�n��Y�e�
�~�,F:"LQJtCG���������ј��D!i�ٞ���:�&�܉.}!�w�>�>���.cn���ׁK����_O�l��o7���X*���8��%���mW��,� s�.��<�n\r%Jϯ�"�hJBQY�l�B
���t���)8V���f���ḻ���{���C{UlMG�M�i���}G�y�)��0�a1U�Y+�ޠ1�б�RA�fd��i8�G��1䘃��7w��i9j�dQ6��aє۟��N;v��?���Fy7�	���Ʒ���E�;v�z�����;n������x�K����--d��	,~��,�g���/�%TO�&9��oe��G�I�i7n.�p�wd��AJq!3���S�6tU�M���hzb����azQ� �7'$���r��qE��џ�����},�e���[�t?# ���W^QS�s:yV)������l��S�Y&��^�Z�7�hXIY�X��u�"��J�P_
n����#�x���'��sTr+������8HE�9�|�5b��$@8/er1c��(��|�qIk���ZW���J�$O�h懓�8iYI��+,m���o�/N�@$u{)��X(�p�b]Z�CG�cs�m��J.[Bx�?��"ק@1����KԈv(���XQ�P�^�W��ϻ��5(��B�Y����i$���E0�����g�*<�EVY�Wϳ�sS�_��3::zT�^#�ǦɅb�;�QjX��%���Qa�D���G���cJ�TF�^���d:�I��P�>�u��̈��U�@��p�෼G�ۅ�P����x��z?�9�2-���T����G�
���b��ʖ��B�k���v����}�@|<Aj|��	��N�s�r+�1z'a���"���m�m���"Z}�&;R ^�� ���B��Š"�s<[�tb��^�B� �>^)=�C䝛� s��p�2Rͫ�i�BT]���xux<HP50�ve�q�%mM[�W�^�Sٽ���h��E	Q�Ά_�ۛ�쫺��L�$�Oz�a��]�y�OInM���L��:{�*7��Ř�㣡0@�����R� a�8�:����])����"YV�f�Q:)0�!����OC;�dG�\J:+U�q�����(�[e���ӣv�!RS[�~��l�K��/$�u�����$$^��(�$�vx����♸�>L��:;��5��p���>����Dw{�I�  aW�e\q��xa+�O�?DKЖ[��l�������-����3�u4��)%��ב-[>�Ŀ��լ���x@6YmM^�fg����ϥ�����_K��d�ypZ�Dqril����j�Q�B��ӊ_��/�typ �2���Ж:�a�:�'0�N}��D�$����c�=�����b����D�6m�Mhj���Y(Q���p�)P }±�7�u�ӗ�5�5�*���X��a�x��h�ۯ�_���%C�Pt����`�"�:E�Ly�跂��"S^�s����͗�	�X�#9H�w(E���ZJ"r�"�F��:�pV=���n
"ݬjN��w���T#��6�8��ٰ��G�K!j��17]�9:�Z�
4��׮��Te�9��������wfbS���J��Xi��'�&n������֗�B�?�ٵ��J�N�'��� pv�j>��̸"��Y
gu��<�R�Ͳ6L('��a��%Y���T9���p�ҦH�O�e=�R�aQq�v�"Za�
���3�m嶘�A��k\��0eO�]b�NÔ���:vh?�e+Υ��i���|M>Ӈ��c��Ē��t�����>�,��q��ocϡ0��[������_��R������,�uf�pַ��|:A0��CA>����Vx�maz�	��x�MD�*H�p>�/����}V�٦X��\�VU����(FcVr�l2nK��@`?n�з6�r�4.d���%�j:�%tR�*ƥ~V�S��D+9�}���g0����{Z�6`�
u��BI<������EÛ��hnR2n�����8�&/C�b�H�(�Q�-����oiM�%T�ky=ۮq��(v@.^Ӥ�:}y �V��.?1���� 9���y�<'X������>���Ÿ��W%��h+�oj��2���ZC�N1[��2���¬� Lልo�U~�c7�h&�o�����B���L,��ن��ٺ���EZ�r�&�;$_��o�2�x�"����y�#�'�mRu�֎懎�@1�𙔺i�On�\�0{���LE/MݯHЍWc�K��
BZ�p���ᏼL���gwt�7��`
��;i��fώ�k��O�jbY
����-Yv�1$Yܐb2�
$H�4~��!O\^7������<ֽ�F�3am�K� D����>�;�ZPm���3�kotE�})>mQ�4nycn$�Q�vU(wh����VAg���?�1OJc
�A�=H;@�u��X�������=��SE�q�Iiۓ;���!�r�*��Ƴ�GM�����ulp�	 	_�4�(R6��(��ǎd@�����mb�U.|5�
mO��󖦚��J"ذ8F 2��z 1�b/b�ŧ���O?z�$$�Us�&{��}�B���ޭ�i\-�5a��s���)D�a���8��!��z��-K�<��-�W��#/�G\#oTbY�����F@��ý�w�8](��7�J0K�ݪ�w��3'{�)ϻ�`�K~��z�Qw��/�� �R4a�駜K{��5r��vM! Z+�p�������ӈM��*=�4�����&�O���:����?��{�������3��<V�Y	�����]Pi�����4�U�Ƈ�LZVtitF�XQ�d�x�`�
��)��<��z�	M�]E��� ��K�"�yA͠s�z����:�b̰���I�i��w�,�dU��j��F�Ϊ��`n7o��^��5�qO� I{��j�i<�F|��@�j{���o�Z_��d�H�Ķ�Y��������k\x�w����K��d�>+���.��vHz]�:�vO�B�H�2����S=*	�T0��3-u�v'����7n�qwY����$ z�ޫg�һ�ݨ)P�;���W�n ir��<u��kT�+��d!�b?<o�`ꗱ�T�p��{���|������E���oL��k��9�-o�hStyeA���LtƦ�P�j}��!/ͺ$-q_��c�IH�C`��i������	�)���iY�f%�����zfQ�F|Y��\FE`�[*��"�E�.�èB�g�2��b���'���cG���`��QBp��mH��>U��2Xp��ǯN�P��n#k��y �d[�3-�iJ:��"Y�4���˂a������g��=����*R����yr]���*Yy`�<`�`7{�� /Hy\�a�Ɵj�Ú�}ָ:Pt)��,�=��L�
?����z,y��gf�~�D5��oofy+1�3�yMӡ���%�Xn�z��ʚ��ˮbh���b�O3h��%^�Sq��	a ��=7(�x&6A�lT5���ٽI��ZBV���H�jͣ�Y�>��AQ \y�P�]���3S�������]��w�R�e�J��A����V?�:�5�rZ����|e�[lk[���q��iGܘ��'��;���2"���P��1����3ĳ@�>��k�,�\��pEk��ф�x q�4NKL��q�/�0)Ց��"�)������/�$�Y�ƴ^=A��z��U���z�}~�q]̡U��d�Y?�)��Hߺ���y({�8��n揤:�tB�_�(�L4$��<�O}�E��{mﯰ��`�y�vv��_Sϖ�`��1>[Z X����\�H�|,��k�'��y���!�6Jv�;�j�l�s-�7KI�XFv�
�u����h9���X�>�+Ϳ'@u�ɢ�UQ���Լ�[�H����#���J_
G�=�DH�]���i#,��k��q�h����gP��I�:��A�62<��&7���BI�Y���A�Vt�P#����bo6�	n�� 4��Q��B&��&������EK="2�W,�~N{����m�A�)R�����0��?�bM�@�|�2h0�o��\�ȑ�A6@oO�`����^��}�����u���w3�x4-b07��Ӝ���e#'�T��gu �*����Zg�_���O~ڐg�j��<�x�q�Ao�����y�j?0���Y�z+�{)8��,��x>(L ��@f>� �:qI./��q�a{�l�>D�:��O#T�P�df�nC�r�]��gI@�&NMv�@�F"q�F ��7~z�i�ɟ`P� �v�n�w;T���)�N�y����#-G��E`�o�+�` ̟�>{4����>�H9l]�A�C�l�&0���Wn�a��'�+�^��iG����F_�g'3����p0�v���j{�f���Q��I�P�i��*HxՒ��hc*����~b+��Q��P~�T���W�&��H`v�4VR7kuҨ`
��{����_gP����&�s��E�}>O=yȲH�4,=�@Q��O�f���������oщ��*#3a�{n�=�sh!;�x��_�C�"*�Ť,�w(Z�T�;�	�2�����oB��#,J��h57��֋�$?:=�F���y0��/T����l�D���"J���67�Hu�[�@�7Q���7��+i(��;r������W�;\4Ү?����CJ��)����jL^+#�v[C�Pfl2��5Pi>,/>�_���B ���R~۾B�p壻��iӸ��5����PR+kQS�n��/Fn�B����1}:��ӈ u/9�K}��?�L*�IB���Uw��Go$��^���̽#�0�ϒ���_l%�#A�g����E�:XaЀ�}��������k�g�r�Kg�VG��5|m�2x!��5��OR�=md:��{���%~�dkH��	�#��[���r�_�ڄD?����l�( 5p.$?�*9ѻ��Ч��Z�����>��veϋb�\v]0[����V��Í�5���=�20�bI13����=B��v�$ߡz������X��ca>���
�Pd?�N�3�u]�s���H�xZSo!��=g�vstz��E�����`�Am��@z3{GE���%h�FM���w�3��+�$<���{�:B���_���@ӡ����U#鏲�3�V�Ԕ�����2�&�r�&7����ѐ���3D}�}!*K[���Kʧ��#�m{6���7��3O�Z��kr��gO{���Q��, 
��y:�7P��Pc�+����45~p����mp�dme�5%[Ce�E�d �gbRa\U}D��bTN�j����R������8|������w�8�j�<[-ǹc7BYO��\�����A>��Z������k�f�\� �I2X���y��.w|�)<��S�������
��!0�E�������R�_��|�W'��� H�2��po�(��x]#/UFʩ��V�̹�"���^�+ Qn���>��{����R�)%�7�֯+X�#��Z0T�U��Y�}�S�"D��a��^$�k�E4�v��~g�у�bS��1���RL�Y��g�ٻ삉wv�0���<m����4�/K�9���J��R�8��94)����Ũ�cu{��~�ә��3���;s��\�%�^L�� ��bWP5��u�Fz
�ǒ�j`�d5U{�F�����O�zg����&�`�9�p�e���j�d�Z���1�cfӟ��p�o�2�>���)i�_�x���X� � ���$uzc\�)!9/F;�jEgqa��@3|�&x9Tvn��f�w�i���	�l����Ҟ�0�Oj���y�M��q���@����I�m~w���Ց'X=Ýf����Z����7�=,��tMѤ�C 9��5%�c���un�)�Fw��}>�����܆��w>���	�8Rd����d��Chq�<~Á@%�<<t��DX<�HI�#���5�>��$.��<ñx�[��龍l�Co:%���*���$ HF���?��Yޕ��K�����x��:L.����ЄL&��7�:�Of%�fM��2rT��@n��)���0
�Tm�����sj�����[#���26�����e�l��q�.G�e�Bȳb$��'
��Nу��n1i���ֺj.���X��$�� ��nsk6L�2��_� 8_h� ���:Y)v@��s��x�JX+ʳo111�v�^�@%�*5���3���p�c��_c���\W��5 qu��s~���'5�e�"��8Π�[�$9��/v�ߠ�ђpw$��H,Ҩ?�Q����ɺ+�>s} ƍ*��E���0ﱈVo�P5Hg���s�:��A�]�:���+f�gg�E�6/G���_��m9!EE�#��/"is^�{�sѶU��e��E��*G7��)`�@EձI�I&M9�(7OF2F�]̣������X�>���c�˾.<Q�[�L),�?d2{�isc��!������*�16�]k�P���̠�cpaq�hƟ6�jb�T���T �fy����f�Pԥ'?�~`nu����%�4��#&>������ЋP�u��X�M*qN�!q>���`��)�ښM��gE���Jg�m�ͫ%i'��p}����:knV��bO��Em%[��4n�+a����>=���H�nKG7�ڪL�h�C�5��o1���b�n�ׂ��TU�=��������(��
��%+�i+&��7��h�a�H�0k潻J{=='�[E7ި
�[X\W���.ǯ|�Ak
�Ǚ��4��������*@ӷ�$%G�$�b�ڜR�t��{�ڄ'
���!�W-@�O��S{���~Ku)D}�-;k�*�m�����Ru3BU�t�c��i���>��U�RCk���h6�w�;|[<�L˾a~sYJ$��P���6��բ�`}x�fS�V�y�Fk�`7+N�g������BN)r�p*� a�{D�����o@�]�172��#�5����z��#yy0U�C��vZ�c�,��*�є�l�ە���n�&�F^�_Zpc�G5�����^	���Y���ɫ�r����FX�)уg��b�ŅL�&r� ������D��H��
�O�H|�e5����WY��T�N�4�ą[a;����?������yE�1��H�Fצ�r���M KA��i˄Ռ\ڕ�Q6j���YR�Y�19��K���hf�b�NYm�Q��/-�����<�C:�iJ\�[H��FB��/�˓��4�����Z����bIQ����eY�Y嬀��<�Kk2 <`*���W�4����l��}~L�K�_Ɠ
]�v���of�#����C�P;5ۂ������u6�!>�?�(ٔ��>w����M��+b����V.�HJۮ��@5q����]�	��qǸ!P��P���[w��� 
��Y�F/�ا�����Z�>��_w���oi#��<{G��&��1)���u��]B�m��	ּ7#A*�-X�U7���V�9u5��y(4v�ă�C��v�\�,Ԕ� �c�W%c���
�-���Љ�3O����Z�|���v��fo.�����>�M�x���&�[y��f��S�M��.�����ZQқ���#5ɹ�Q.����-[��� a��Q��5��#�#@_��O��,=d�j=��'��oƺ��Q/\j�O� �{"�D�2����/��׃-�����Vb�7�pV�fv"
�-�ܑ�[���ZS��jҷ</7wGñ��2�Z_ RbN����cK-��t,-*�) �ӻg��jMv}R���J^=�]�ɔ8Z�d�
����\��R*�Z"7U+B���If�U�f�{c�C�{����Q���@��;��
T2�l���*T��]��a���ތ������JᑬPB@v�z2f�¼̆�R�м��V�}L��q�5��ٺ�F����<,[���E�=��	n�"ˡ"�������( �K��G��C�幥��m����"�����9!��|1ȑYf#��Li���*��<6�V��H}�Hӻ6mj-�§��jBl9�Yԉ��k8ܡ��ы4Us<_v�%đI���R�����AG��-LAY��V��zŭ�3\����þ�m$��{�����z�e:#�+4v�~��[�m��!��;'9� zp�΃����#;�e��U���c��uP��g	�LC5Q�-��]��jp�Wvg�I�U�9u��ï��z+5k�ut����1uu�půs2��^����DX��aUڼ�ld�鬧WҨaE �G��x��������TQ��1F��{H"���4���+�o�P�������/!�'�o-�Q�
M�FT~�}�y��sU���8��(f��`�."a[�t[j��������T5w8+i�U��]{4��Y��ƾ_vi���? z�u���׶��_���M�ҋE0��x�oN�/��>�� 7:����� ���׈p=l�����΀*g[+��(μ�.���7�:�N�s��}�����V�A\�֓��jd�pgVV�����a����=JCs��Q�sf0��Q��#Ì�?~%���+���3;���}<�����tM�cy����A<$	_��xgu�z�^�*TPϲ�Ok��&�l���>ͷQH���Y?�d��v�}r3܍Bh�>
��+i�/&��	��Z�<��\�?w�X]t([�8��`����Qlf�)�f�3�B��#ic������n�on�(7g�*�G;?<�whqGJ$Ǫ�qY
���<����N��)G��{׼{~D'+W�΀��
��󀟆ktu5im%��Wb�]-�۬�֟?��/%֓����Ê	� ���7���i���2�u�[P����j%Q5&;�J5�HJ�-<�a�|����'5��cr-]Gz�B�X����hX��!�A�7�%��H�J֥���c'p
����Tpb���M_�[!h`5�O�f�MF�]t����|���]���ӳ��c�K���z�^�~w�I'��K���c����J��):������Xz�	�����6!�?�M��6t�w��-3��I!v~�v2�s!x�/�+2�����3�g��i���%��;���W��"/ !Ժ����3Z\W�E g�w;6��bJƖ���O0q��T�jo/�!������Hn�j�+���/�V��k$���f��y ����<Kq�Y��.�j"����t��L2���4+S��|=jo������D���?t��N]?�V tZ���n���Y�&<\�|��'j�����4YYh�(|�3� x$��P�����
1J�x����qJ�FN�fH���rt�@�\>di+�A=�G�Z�_�x�_�UM���/��QI�� �;,�UVn�Jc?�l0/{�r��Y8kx�mt�Z�6�)�>�z��+H��M��S���}=sŲ�,]>�m�kkk��`��VW��y�Q��1��6��H"���	W/��hn6��ΐͥ�
|�.��,|�\K��z?���b���8W�ҶPp��U�������RH��\2�b'�����Wj���*�Ԉ`��Sx��������f��(.k��yb.d��尮��6�q*�,�yK�_HM;��K�qo�sߵ#��@��R�M#��Q�?�uҨ�����ed�Z��C���p�aYA{�m9��B�F�Q}����o�hը����'�����>�	��1�٥�JC�cXQۚ0��ѻ���x��T\�H�� oX��N����S��?%��UT*�㭕#�q�����jꜬ>n5��mO����Y5L�v�@êjj?&V�|ˬ�[�������1U.��q0�O~�Sᡭ��z<n�����`"�����t���gЈ����Ua!|�x^��7i����8>�,����y�vA9P@�z�׬$�j*�
��D�H�����&�~�l�|V��@�~㿄�[�`��O<�(�d�߲�Dv]F��P
��B��7�zX�,������a1K`
_�����4�u���N���ԝc���K}�,r���~u���p��,�}�e ��o]85;�Ĕ�"�@�K��bK�ɡ�죸�e���N�|�J�3n��r�`R�صnmc�iW688t�kCOO=[�u�2��p�x�K�؇��|\62Yl�O���0����]�fjʯ��󦿘`hX�~��G�p5�i4�]=�:��
������:F�^?�fNn�t�pIG"ǹ�>,vo����a��?>�[����5�PJ��Ћ\}S�����	FE��cZ�s�[(b:-lG��]�艠#��/񷜁9tX`,��?���>�4�i%Y� h> 1ZY��B1Mݥ��R��v:�8SR��F��Y�~0���mۨ`@>Z�ٙ�s�<񭭩�?�J��m� ���gve{]���i��ͼ߻������q)V�5�A���#l�}s��"�W�`��s��,l�;�c ����]�kdK�k�ǎ�.!�;���\�hX�8�/��6^^
�eg瞮�2���S���c�E�s��JM�KAHX��߰αc�ﾵ�{۴�&�jc��b]�Kɤ��9k�R>�$�k#���+����#M LJ�����ƞ����V8tc���A͖�>t�h����#Y����k�xl����v�w�����Y����ް��s����;��R��'[��䥜�k��X���/��r�]�ģ������^���`)�	�VA��Yֲ��׳
�߭z}��}/�bh��W�,y����VS��k�eD�����o�7[/,	A��n3�NO�9��ïBWy����G����Ѧ0<s��(P��Hp3��X�\��`�L���A��J����`%%H��-����|���]��[�粨ۃ��vL�<�1Ʒ�L�6��?̵W,��I)H�\7���<_���0\üԥ��ɝ�k�S�E�.p_۹V�t�C�΍}��#WC;��']W/pN�5 ��#�Շ&��cgd���`�7n��4�����4���>�
��i����v�y�<�]E�y�^�x���B��~���GT>k�cV�06�~j�s���ŴlP>�Ý;[Ŋ,��"�C�g�.{�~\ы�(�%01ݥ�T7���������ū+s�g��p,b�rҠ�����_	QF�{�1���&n��6�I1¸b��������, �f0��S�_S�&�:�1�;VwP��^�@�ha��C�q	9���t�������F�&���},��u�C�n²�R�t��OPY�U�U���K��;v�?TM2����y�Pw}������-������,¹	v�rɫ��)�@����K���^��i3Z��A��v3ͭ��}�C�o���k���k���4X���뫮#'���1W�5�x6�� ��ܼ�����˓m�e�PF�����z��ʍ$��7��KJ>-#��=��i�K�5���ԡ� `n��K���k��B7�K�KK0���b}��T}\��7�6��-c���pw���e�� �?Z<����5Pn#~|����vM~݌��gS�`�Y�8��\Mn�=gZ�aչ�RZV�T�D�#������7�x�0�F��wv���N}N|\�t�י)�o�w�9��cc�I�_���c���_���x��8u��6������^�S�98�"D�nQm�E:\���{i��|��O�^g�~)J�S��r�K!�=���S��m�K�8?[�G�/��:�E��`>����>0�� ~��A���L˟��T�>:#lI��D��l��ͺ�1��諔#e7F~<>Gx�-#~�Rד'4�R�:4F���̓�Ca�;C�^�~E<�2m1�����h'�Ӯ�T�o<�Ɠ�[�D?0`SU��Y�n�Qz~?���4c+*ԡ���A�ǃ�h�Ɠ������}�q�hR0t/%�!�������i@ּ�>;��}��V7+	��ƚ������w<,�����Kg64�a�`R��Y{S�������wR�'+�[�'�`��et��*-̍�咱�����?��D^�(V���v��3H�z��2�T8Rs|��"�:���ˁ�kg?�D����?����{���O�X�#89�M��Ժ��WU�G���T8��� <�+�,X�'��ݮ�[�+r�K�A|�N�>y �U{χ�Z��_�2�h���k0��O���/<aDS�U���������Z�lJ��ol͏�m�U���V��Vmɳ;�����pA��m��P�/j@:_�'so��g���54��H�ռ�F���nJ��<wO_�/Vgˠ�a��.��J�[2�ZY�l-�h ��
���V�
�32���T��$��M�w�G�`�z   �ݭ���f�7��&�qz���r��/6���я:򃞃�hk��g����NNm;J時�Nt��Rn����Ϳ�*�"7���"�"N�0��s�,�LG��V���/-ۨ&�'~>�;����R�Q��H{bIN���� �mG�f���*[�R�5�Z���K��i��!z��b+e��;o��x������$$��0�)t^���4��_��+-[z�5��VS�wW��ʑ���x]�;��2�@L�D�?R�����*e|yrg\E)�x��)��DV����������bP�p1�����U0�N�����q�̕���ʷ���0��G���F"Q��^7�a0�^@t���%��[�ԽN�<s��	kߨ�j�J���dM�S�����d"9�����Y*n m������l���Gg/��mZ�f�6|����N�p)hƥ���z���+V��~s�t�	02��h����FX(gŗ[��Ġ�Z����Ɇ���F�(+�H������I���/��e;JԘ�V}T�q{���(��e�g~\BO�6����(:�n�k6��e���99��}��.���Ҥ�%��[1�jo8 s�	�����f�ry-t'=P�H0����H��9u�,��IH��F��tcN�?j����*�������S��-��'�����3x~~~���у�(�8��0���z��;p�k)����D%}y�����}\}���T��E���h��#:�A��r�����UN��[R�}�x{�=���,,~N�@
�S�iwZX"�?][��$�u���ꕘ���u{�y��{��|N���X����qm}��Y7+r�UQ��QjX8�՘��{���5;6�`\�B#�`��T9$]�O��Q�LB�ԩ�T]x01>�vR@����UyI��P��O���o�
.�k�P4�}�E�eW��̬���77����wO��UG���h-�oW��X%�L��!P����{�5�^w庻%{;=���|}MF��7WLJ���:cW�|X�8����w�糪���]r���;��6�Ѽl)"o���,.Vy��P�z� I�2Q�E|aJ��rh�jGW�A�&q��.ǈ%��T�P��.�|x�g=%������^ڒ����lQ� O��m���%P҄,����||�XG�w8����<��\[��۲4-f��<���@�>��c��Ѷ�C#*t��$�O�w�6��]��K�ђ�s~�fW;q)3��>�C�Y�����A-�Ǜ�S��>V����j�9���
#N����&�d�n_�7��6|�$��;��*ka<�/� �g�D���ڏb�\�/`u�v>�O�15�����k��;v%� �c���{d�d�9���c�_H��6Qp�\���p��kx>X���5G�k4Nm�P`�E�Tt8�^��O|���ީE-,:<gHB�'5��Q$I�I��6&��O{��ׁK;0��$�ޒ��!�;�(�^kZ����Ky�Z��N�jhOn���J\�G0�!O5�����y!��������E�ꀢwS���&�o�>̓�17�l�_�[�](�
�"_�ʢ>��cϊ�C��À!�	zy��8c{\�"Y�,���#"����o���}�֒��+t%��H��o�4(��?K~G
��-@�?��rG�Z����P4=�'��ܰ ��û���`��Kp&�2Z�T����X*��-v����=-��
���g�'������䨰lה�)]�MN�K�"��A[�{��.�|����4C����b���%JTY[[j�>��S-�Z[�>V�b�18�=w6QA	,`?:�f�֯pm���#�+�.�FO7�Y����T�V��O����r�l���Ӱ��2�$l��.Շng�]|�z\�W�2K��?1=�[�BK���������:�quq�c6���ʨ��IByyC�wq���z@�wp�/ZIi��N���:���.SUE��Q?w��5:��\�����;Hh8:܃�HPsE	�o����]���_]}���I(��*J%��5P�ꕾ�:kk��JsZL�l��y�4WS,N��66p	��
MO�y�L�� ˶x��~=:�5:ܴ��h�vw�
��u��W�X�T��V����u@�W)��/=k��N�����TR:虓�P�i9������|�/�ˠ}�7�Ι��U`�1�&�����b�h{B����Q論�_��=q5�����Gj���*V�;e��ȹ��Ζ��dkZQx�oҴg����M�>������+� k�v��њ0cK����*�x������ǆ��{wq��w��s��4�ͥN��pxe��w8�k?������@�{ۓ	g4˻`�s(Ԇ@sҘ�\����l�>`0Z1x��������b]i��۴^�'����it�jV��\�rs`��\�Bu���m�	mL��f*��=7���[5s��]۵����i��������.q��)�ˎz(<��`h���P��O�o�s��'Iʰ�����w�ؽ���x@�ۤ�O�>ͷ\���wc ��2ld��?��S�˖�1 �?��W|��j�|h�m��^>.NʊU��W�0�v�ua�p���X忨�A�U��^c%�[��&�߅z1���xJ��9Ƹ�y�����RCS̴���V �߷����2��k�� e�tW���MgU�~�!Ei%��E���A��[���A�[$�F����F����=���χ��쳯k���{�;߫,�2����H۝5��7Z��Y�VF7��^�k���+�B��x҆O�R���LWr����IG���;,�Ŝ(�?,�Ṉ��~ޖbtr�}��󇏱��=�
{�ҲC y�Y���a�Kt�[��@?O^>$��x��\��V�����7���=ϳ���*�W@|H��zz'Wm��4��P������܌��|�Pd:a~�]v��M�VI��$���^s�i�X"58��xzz� M�	�����=�v�=��n?~�����C���q��/=�K_O����hr�s��}�B������U���59攢򭖓7��mc�f�m4L^j�-����j�jJ�8o}=1� ��wv6�g��c��G��|�e]��SD1H��y��V�H/x�bDc��t]ʿ3i5��vC���&T�y�C��5N �)��QI
��C���DY����@�o3ޥi�$�/^���4����z1@��V2���jb���i���������i�/��ތִ��̧�s��ܾJ��#,
�I��n�9�����2 ]ѿ�Ж�߈����G.��x&�j������ROk���6ZVx�#�=� 7�:�&�*Z���)U���R��Lmd�]9ڢϑ��d�X?�z�e5��-����	��E�iY�z�����s��q�>ŬvY722G���k�+ú����:F�:�pd��p|����Aj;,���m�ڇ.g5�Jļ&K��0���v��H���V@5��T�J%B�"u������golile%'���ϥp�7��s���=��iY��8����#�p:���L"_�=C���s�^Q_�.�;~D�!�|LY���n��U�&�
�a�1��6��!]�ߙ/]'��hS�����������_Dy�5P`�j`����N�8X�UM�z"�{U�5�p�,8�.I�L��_���߿��q�Ve�EO�O�KT��&W��������x��'%�����K&���	�o��D��%k�>8v3@�pU�l��d�
L�LGߏsJ�k���<c��R���z�4����l����k�=O˟��.u��|�8|l_ڈӯ�bp����J����ݿ[�ؙ��ݥg��"+tm��k�m��A3��]l3��~.�����~~v�S,���~�8u�;\O�j��X?�	W�5$���o��S���~�V�����ݲ�m�2B���d.56iG�m�\e<�D/ � ?@v��
���K��g�E���R��i�}p���0}�7/�O�g�N�$���5�����Q���H��ʩ����_� |�]"NQ@�1�!y7�n�ka߀7�KN;��1-�G8Gd����!��罓���,�����\��X�br�#��!�N1�h��\�m��q'��&�A����g. ��LF2b%�%3_�F{�F��a�����v&� �V�tU���I��F�fy��6z�L���(���og��lZ��AC��0C��0�+�ZN�~�s�¬s=�_w��pR֕�d>S�t���nS�����}��`����4Q� vN�6\��.��"$VւcU	ls~�^��Ĩ�l�F����	�����C���y�s�?c��v�߯=����,+��s޴�<4~��N��B���iF������+S슊}���1�gנ�� e�UWg?���.r؎�-��������aݏ�$��wD�{z�+�:�+��d	���G����p�`�"ȼ���P���ʭ��䎳���AhX�o���kŻ:7�(��I�<H8��	�@;��w�`D�	y�i�Z�F2{ڤ�tv�O�Q��o��p3�Ou4c�w����1h��m%�k���������㜇�LbD�eC�����ȶ�b���XIp���������9Ek�߂Q%�����u�1V�}�����A�">Ԋ��]�l�G"�Ӡ� ~)�myo�9+P�~�!��Z�̴�n�X?~Nz�O��_�֥�S��ʡ�����+��7�|�ꑙ�rƌ�]�ٮ��}���߃�{qN��Jr��T�^Z�Bw^T�N/A}�L��:/��X{��0�q�;�����������
2���:����T�ɬ�J�\z�0E����w��\]�a1�E,�C�62���Svk����d/�7i!��B���ʎ�<k5.}�?t;6��<�m���SL��5 ����;�:�G&��W�G�j�G`#����|��U��{^��TB��0)���&k�����mz$�N�Z�I�0hm�����AE��5�8x{�@�֝},Ϡ�R@�Kr����^���������I��sJ,��NayAԝ��Bqz2	?�� ɯ�B���e�t�ڿm�34Oɢ�P)q�Ęg]�0����u�ߧF��9��Wn�i��?��и���>֗�\���v�ױ1�������[��wd��ԟ�_~���s^"�ܷ�:an����{߸��K%:4̜kxo>�f�*S��t�g���1�(��b>�鿚*C�0sٺ.dG�丠]H�С{{�QXh��v����i�y���*�6����MC~��=�/B����.3�o8����&�c��2L�ֿ�Dd�6�`�4!+���jk� ������mqp�XG���*��}i�d�Bɑ���ς�����_c�h���dwW�-���Ps����e�|���'���P'��jV�>�'�6�C9}[��4$�1�9p,Aԫ��{7"�-�]4�I�Ƽ�B-��@��+8-2�����l�|Rd*�H��֥�L@u�á�#3�Mgݖ���_��T�JĦ���¢:��l��4�i]6~Ѻ:�����˟k޽�ʣ�8K�%~�}��;��Ct�|����#�VY�VxT��Uf�e-3ֿ`{)��2�#n�؆X�WV��5�>|�\�-=�0bՀ�ҞAQ�A�9�7ϧ�(�2���d�I���J���L��ǈ�<���l+?�QQ5���5JV���RS�aJ��{���VZ���[};ˠ-�b:c镊&���z,�0���\��ǣ�є�sYh��֛�����_����c䨬������R�>���۝벗�?h3�F���[+SŞ����rh���	��a�)H���I)x/��L���2�"?�A-6n��m��A���T	�2����Q�	��vދ�@�}���l�B�+7�w::+g[�չ��{k��i ��+�DC}�f��V�-��۫Ӏ1�|*?*!��sa��FP���3��U&�����`��&%e�mGr��[�m[+w���2����!��G�>k�t!$١H�����J��k�q��>,�W{ONk<<:zlD2�_�ONz<���Q�Eg�l�JsO�[MÎL%b��	�߰����b}WE�6�y��_ف#�� c�k7�qm�=���I�\�tG�[�����\l�����ȱ���f�V�S����!gக�Q[���)uЪ.��2f��9_�#i�^ tJ:LQ�_�z~�z�'-�=���vQ�a�xRXR^���	����shR�)�'kJ�Zs��l[�[�V]�B�1益q��f��Y���c'�.B�qK�q�����@�~��!��DEE��}^}
R>3�yCX��j �V$�;62|[�}�1^�N/C�dVOZn�;Z���lT�I�R�~�?௩YA=� ֨;b�T�΋:��V;$��a���x�j�c���k���p ��<A^�S0zCO���ο h�:�@�Fq懚�H򞪗7Q(���S�������T^j�>����D;�̊���b��0��Jl�������]><���ׯuUK�D��Aĝxhp��ߪ! tԉ}�+߻Rj��j0&�Zl��;]!��5���m��^�L?2���}rv�:U��3�Ώ?�t9�!2�Z��(\����c�Y7�uJ|�)�$cha��)n[�I@}�"9x�����4�}J���Ҳw� i�DD|�󞙆a�'%!q�A��Q/�G�1�sko�.�ϋ�v�C_��O��]H�tSUQ���nd�Sz/gm�Ĵ^�sl5������.'��塢$,�N�K���\rg�3��^ȝS���Qm�&[�$s7����7��p�8����JKqj�����I��b��󬵋T�l׋�n��7�^��%Ϭ7%��ht�Rʕg{{�|��|bb���s&*>�.N�b}���#Y81F�D��3<�)+�K4k\�ݴd��cK��-��ap��@%���Gy�� ������m@5����Z����-Ό�"��~�Y��c7D���ZG�x�W;c���ks%�ԖhE������D��"oCV���#y�V���C�B����a@��C(�CD$1\�c'Aȶ%7yu�'Χx$n�6��f��OF757˫��
�6�U��w���n�cm�u�v����-�J>�ɶ��[���蟲���s���C��H{��;���)�K�7��f�ұ��@-\j���a������D���p�����[����
*��ʸ��@�+rr}��t�b��z���Z�X��Y:��>�q�k���_����ҫ�fC!�'�ɯ��LfZ#��1q("Ex��� �tw~�Ŕtc` �4�T���o:cd=�9�Ix-������7�Lx���o众"�Lx��gT.wVt���i�o4�^f�����2�fY>�5Qri����O)3"aI�����!2�K��4��O�!9',�`�ۘ�B;>~(����W�Z��X��g�:����N�+=��	_('����u�_�r�����*�q0��j�N�l���L[M¸�Xdx!�W��i��X����1�xZD�T�}ڔt�����Z�a��['�#"zt9a�1����wO����_��������<`hQ��*q!�	�P�uz���A�	���(��W2��˱�DJ�9Jbz�6A6�.��7A�|i/�SK��$�/VV!M=��ڦ8��[��聳8��/�s�4nwW��f��A�X�l�GVm���<G�UC�`��"�1J䎜`��^������E������s�%r��݃�c������}*A����y��ᱵW�匛���8�=���M��[4�bB��O�f�v�ȸ��X����=LB���;�"E�<���M��Q��2��3K��,"Da���ת�p��.�����1�f}���TC�>:�uu9��s����2}������սo�0�#BEO�A��_/�
e๸�ʗ��S�a�ɜ�O8�VGA������X~������_��e��yWKF���a^�j��i����>��d�݇2An�&��6&/U�����7b��$�x�(�B]v։�tE&�z܄a��є%�fk��8P����M�{{/�S��z2%����u�mݙZ��9>��������!^�/�tGh$�;���W(nK:����4��cf���Ϩhu�����Zs�w߼����We&�$u9�{�~?��?�y�;(RvͻQ&���Ġ*��B2���T� ׼~R����CjF��DRa�1�����<� �C����.�v>�eOF�l��9rˤZ����1�eETux;������m}��[�y"��e,�j\4��HR�Ϙ3UV˕������7����FF*��?��,Ty��eX�6�ݹ���r�x�-^h���EK]��	{g�4�Xa��@
��`����g9��HG��\�рئ����w��CO �c����&��?���جY�t=�W&�m�����)Lm��\���2��^��Cȓ��w���BB �#C�m_�NLA|Iu�YmXK��z��e��o�[E���$%��0J#[�=�ga���z]_�:�N��S�K!�B��a3���MI(����o���}�����3�G�d%2�S���.9�/�T~Y$�$a�3x��HVL���Ցjn|���������ֽC3��҇�t9�LTP�4���J9'�:\��] ^��p�U�\�h)u��,�����5�"Gw��Y�cs��,y�W���SD�(�BW'��|�v�uǋ/&�}W &}_3=I��3ܖ���؃6�fe���V�Lk��_�@�a��Y�Ư致ȉ��������kyE���^�S�3a��>lz|�5Ж���]�������^̓fc����Ek�'��� ��G["��@�C�|����_kr�&aP��Eo�ŷc�q�[��;i���>46�H���RsW�<aէ\H��4��R���5��ūF����˹����끶���N20�>���s�����KA
�0���7�f_�`�	�z�Y����O
�?w�6 ��q� �~��}F��� 7�k�����Ŕ���Zc�~Ԝ�f[_z��tjH@8�]uo����V5����m���́~��y�&������w7TbOL�*y]x�=�'��SVl�U���ܸG��Q�I�,Y!]F�e\T��m8	���S呈/��^9�9[�1'��)A�Q�qDs���~p{���b�, ���RiȠ���؈:�=�3'��U���'�y���'|nO��r��7��,	yZk����ڟ���1�$;P��������~������"��PB��c^R)�إ�J0G��̰�5��x~�=�Z��+P���?�t���������K1%��Y���f[ķ�Kp{\����o�����7�4��y�H��^[h��\[uINX�w'���kC�ܩ�8Y����;�f>\V�wg_�F���)-�J�+Æ����iR�Kݟrn�~u�2/�������rg�L�k2ѳ�v��4�]�����������v7i�f���=�+Q�F�ë`�38�N�͠�r�e_��nM��\\\��7b�U� v�w�8�<5��zx�{wC	���2'�-�Q����o|M�r�s:"{�����M�v~CCCe�y�s�L� 1?��2l|����i���L���������A��2�����2��4�k��/����a,�F�����̣/���)c���]��^>M�t��Mܶ8�*���v�&=#���_w� 8bg5C&dR��������z8<�k��� �(n�hwo/gL�����8�o ��z�#����b[YY�06�͵�ѻ.�cS��=rZ�SY?��^	��&k4�\�斾��������H[��YC�@8j��=������:
f��s���U$/T@���lU%$L��Ю�&�%w�S	���a}�~BO�S�Тk��b�5gв~n`�Jab:���V��lsNG���ѯ��y<i
G��t��@�I#�4JxTh��+v�gg�+�KI�(���QS�^ۃZ����@!I�b�h������f}��3�1#iD�����\�:��8\�pBZ:�,V�d�v�����ڑ�}����2���Җ���t�O7��w��鶻6L�8�A�A���;�],`�~ΐJ��Pt����������i����^v �)f�y��(� �;��F�UL�ٷ^3����}o���	�(V��4wtT6�8aV�.��,���v��������Z��\Z�{e'���L*p�K��T4��(��b�������ƖS�� ��B���W��A�YBrZ~��Ď<{���)Vl�{�~���a���D�"�+m�s��n�@;��%��%?}��x�čLZ���I����&!^�L����O�XΧ���D������M#�/�
�IC��3~$�P��|��� K"��m�3ڶe6�8��[FȒ.�Mn�~�vsw���;�s9��O#�U0A.�c\Rw�/�!i�#�7�=���i�pp���Z@Kd ��4��4��gzi!�bg��u�9୞>�f*�˳q���U����mq@��q��	��?�fe)8KxKgQ�3k���鼃#})��	��-`���m]v�̤�d&}h^wy烑�ߔ�Y�Pa&I�23�-����wjl�)u��L����D������c�f��m�О��,�=M��47}!������=�=/'�������M�ƅ�Z��D+}�r�e�gq��
G�٨5��:��a-ψ>-nd(R$�|xI����=�Y?k�1�\27[��8P��_�����h�}�(;nB*� !���N�lh[c��O�U�q�I\-N^�V m#�DU�>�UD8۟�q��0�w�8���2J�����
�$�/���<�7s�6����N
�jJ�WNl-ez*.��y?l=��F�i�=�7Gtv���<�tWc�ت��--z���,yF)C�2�Ӂ����͊�@�$1?����A-`x!oѲ����8	��/jf�)�w�g���p!֞����ڡ>d��� 	*=
�}�!w��0x���:�_����+G��lEx��~M����egaꐉ��p<h������+�	ny%�n�0��w����l��Չ�[��q�
%ыϓ��+��J+I7�E�"�e9n��h*�o���>���e��f�����3��*F&��7�X��0mƴ"C%OD�"&	�'(Q�`�,�mN�ۭE�ׂ��ܹT� k=��ç��&^�`c�ڋ�Z�r�K�H�h��Z�1�RY���eR�!�3��k��v��j1˅�R����%/��)����6��Y�b�=��K���W�y��؜���$@n�;��iŇß��KoL�_��ˊ�?����7ܚ)HIKS�Ho>�BWS�^����쿇/N�'�<:}i�5W�~w�������]E �x��$+o⺝�F�Qpr͙��(�=��T��&�`������P#���uĞ=��d�1�����No������v�[��ZUX�~h�������k�� Ik����f��<�Т��9�k�����Z���t-	�dgA*��㬮4[z�� Ő�f.��k'g<���,�V}:$��B:yp&oǧ�V������VZ�h�8y=~��/qSաW����k��H-97��2vSʪ����{�v����CCٕ&	����SN ����k�,���l��WF?����1�N��Y���e��a�b"�)��O�Ɨo���������)���;	LH�1�+��A������BЎ}��b'�v]�>B�u�),�xI���l����㻻�oT�W'��э��yx�����f�J�h/}*�ׁ�����ɥ=�P�%�4��@LH��	��F�S2k�-o#1a�@1md���� q��OY�vF�_B
'@:�W"7�+���a����W��]O�ܞYܿ����z�ក�'>��;���!#�d�ћ(v`��X����%��!�Q-=������S�B7F���b_P	�`������&�x)T�����Q�QU�6��/�7�\^֎#��Z���h�\�=�1'q����.�<}A��s���;{D@U��:��əv��o����a<��i���S1]˯��H �X����+���KƊ�qc�I�Je�u��Z37=#�x���k�P����R�z�Ȥ%�Q�f����yᡛR���!G#��T4w��tD�?�������.o����/Þ�}�x�ě�&��{]E�a�Xt[fr:�Dq��eUf���.�����C"r݃��V���u�Qn��鴄�.����.�AZ���q�9� �i z�Oj����$�.YI'e�ǋ��ӝ_-�ɗ��}��	�l�Pd�}"/8�u|a�в�dZ���r<q'���n-S�z�'�����e۝k�~�ʹ][�������뉬�a;/��ƍΠ�PI;w��>ǭ��12c�q��J�^9,I��y�c;hׁF��OLW�����L�\���)sa��-��E
���]��7@�JY�ښ۰� <�1y�c�K�0�H <��h���t�7B��7U��n�Ϩ�@����i��0��g��N�>F��~�8��O=����I΁XnY ��.��\>κ�\�M�I�.��CM�e$8���g�=�"�7[bo�U���� �\�@k9��%�Ñ+�[6�&�{3Ҝ)�@�֎���`�����;}30���{x�sܨ��ҠQt�jta��&����cO:±'3���%���@O�s􆧐�p0��Oj���yX��F>��&c��'������E�0n!p,��+�qx����ȫ�D��\׭q����ߒ��-���ȱ�tp3:Q��o�!N���Z�Q�o�Z��Zp.Կ&�S�J��*�A����e��b����H^�r��Q3�8.S��A	Kb��?��y<��{�\W�D򒢓�h���g�' {�v+���=�ITa�����Q��&::А�뜂�2����O�+���z�Y'��Ǎ��G%�P̿�&�����2�u>�����{_��fs�'�ڮ�^�KT���?�ta��ׄBe��MD��%sJ�2���߶�ʖ��7�	ATJqqBC}�b�
{�BI_k��،�W�%�F���D���IO4na��7��9�Ҟ5�t�Q+.����"�W	!}#�gz0]A�X~䧉�`2���� �泀b�]E��qg�E�;��3K����P�l�%1G�n|u��)Y�>���B�-����{P�8��������Z{�n�VV��.�dJ1T�'�8(=�i�|Ϸ�cN48��CG�H�!*
�z,�u��L�u=!�����*�b��'��ɑ�]�.�&����*3�(�i�A%s{t�����uW�P�;�_��$
�HeM|��J2�TQ �?���ԕ�}��!��?�~�6�Ϸ5��x"���ɬ��!�if.Ш���I�����
?	˹�u�����`��t�Χ�Oy�c$uI�F76�@�oM����%Z���}��U�$44xҚ�(�Ç���zߝ��÷��`��LY^��ȳW��=|K���V�L�jFvw)������?.������+�������s�g��Xh��4�7�ōr9�� q���p�d�* Vh��kZ������Ϧ�y�P��76�ttj^�� U�6��a4�x~h��A�3)'��X�<	/c3�q���3�t둇�u��Mb�5\����X�6?�$*($47�+�9k����=w��6v��գduBB*����s_����7�G\�ZO�����z^7;�(�um]��7N�ַȔ�j�I�~w��!���~k<\��LR�j��F�O������'X�[`<U�1�8<G2�Ϩ�F���J	��
�]�5*	p�WKOW�R)���gԉu���6�hi��T�˕�����Ɇ�@oP@S���8�f&��8�Y
n�d������
}p�b����|̪~\��^0���$Y���cϕ0�����c�#M�Ӥ�E����`��Czq��������žag�����	|�g��s0�^�v�l�7����p$^���
�,9#<nJ��}i�a"}���0��ރOpٖ�L:�2T���	����h3��U��$kG\B�a \�{ X%�G6��mz�s�(@p<�|�X�; #�_z�����������i���H��ԭ-��<M��0.7�����FwLt���tt�e���JwkJ���m8���<�e��iK�����P����r=RB܎=�Ƃ�-C�ĻR
�C##,SNm}�'�[H�����/���%�xӸ�3e
-R�\V�:.�D�3*\U��B7aG�I/��\�h�8�0گ ^��aN�v�4(��qA\T�S�=�V�i�( P\��:�{_m>J����_��������Q��o皽n�y����o/�a�..S��KA
ϗ�I-0r�h �����~=Ka߿ĜB ��#�~�ׇ�.x�-�N�� �^�9�Ns�+&9��>�)/ %����.US���Z�xFt'Z{�/�Ʒ�)Q~\��z��XX{pl[?c���\Xw��dw$�~5�Tщ$�:F�w׻-����`��	À����qF~/���W).�P�c{������H	7���M,���!����f��]���P*�+/�����\8@/��m||�RR�c��vw��j0�((��<:��^ȴ�l���k����\Au�Ѣ�B�l~��A�e��]�ǐ(�ӏ\t�v��	�x���6k��$g(�VNZ��Q�v�X��s���<���1GϪ q\V\@�,�>���Q <�[!�����Jhn�`�B.z��h�D�d����: iI���~�/͍߅�X�v���6��;	t���M>)�տ�8�Q�)fG�8�ȝ���	7L��L����Y֥:L�$�f�jTd��ΪC�@2ɘr^A5>J	��5�&��|x�c�K=x�%h�ˎ��kGK����>��m����V�+}E'��[�{��.^�� �Z�?���)�����s�|pĹ�/�:�om������l|�BăD��t�N�勍�(�g�'����J2��0�F}�2��+�[��T�BȪ.�s�����0e���� y��~�4��%��i{/[EP��� %���6mq�.iDmGF>��0%^�2,gn�#������8E�`��ꚃ���Йw�4�̒m���T4�ޕ��++�BY������9����	�`�p�<�{���N�́�/��D��^�_ܑ7�s����Cʷ�ť�;�p]#I
��9��a����Ŀ��l�#D�Q�9�4K����&�Ƕ�r<�r�S��?!��{�{+?g�v���Q���E�~��Y�����R�"S@��('I�f��ﭽt3Y	�p1�C8dV���ez�6��o�E֎�<���0%��-z�*�[�N�]�d��^�.��f����u� ���r�����U�ڧ=�3!����zb��Ei:������U�L/,tV�z#� M��LA�-�]D/|Z��A���>�-�#3a���kw�CL�f[s5X��o��y�*K� }�͍��a�]'�����%�/޼�"CS�Y\��h���+���Γ�o�\]��\��wS5x@ 0圯�Lu�&�=�}+M��{p�X�%�p}C�vF�e�_Z�柗5Lӂ�7���U?Bڰ��� ���mIr��~J�������m(-��
��L�PZx)#�k�Ee�������nc�e޴��o|U Ot�/���'��N&lqNLL�Q����:uW��hc4��������i$�~�=\��v]~;��?tʃ'
�VA�@�����V�܆�l*��V:m�����$�]\����6�ŋW���>IR2�n�!]�^ihJZZ�Ėzhy��BJJ���)g�_~t�@O�Aoqz5�79H�H�n\@c��Ln;��[h�Q��B��N���6���A|����-�FX���d�g�^�����ǹ���@%F�B�O������i��N����;����WCC��	��f��2M<�|M:��)*gOo/�5��������^��{zF<��im�V+T\�	2��:�/�<��2����x���LgOV��aj��i���j��1/~�[xw���M��#�yFF*��}���i���y����X���~P硇� ϣΗ_����nȗ���Q9ݐ�����P*C���=#Ԝᖺ�b(��:� ti�rMٮ�y!�����w�ru�GA�%��݄�c �F��ͻ�º��� 
k��X~QE�}�˰'�I�\��¡�i*�J
�U5c?á�5*?�� T=KN�J����}N1O����ϟ�?,�ߟ����
^__�F����*-]-���5�M���z��jЈy��DsU�����+�������"L����6C;IC����m����5�PpGDX���(I�ۺ��%H6�3�,933��by�|������#t}�H�%�*K�y���`F�D� h�hTH�:�G�K4��ꭄi���5�4?�* �T�Lh^��0��[�ҥR��t��S�?6>zB �9Q�T?e��>@�GXn߬���G���ԫ�LpK䪘r
ss�BkcLz�^��c�E�W�U�W}��*�r��J�W*O���V�}_sxU���󦠚����	Um��@lg�)Q�i\֍�g�T�w�ݍ�/
�ۚ��G�ݬ��bG����j�A�h�W����#����~[n����d��#gf�S]�QrI f��M�ɧc�Q(��13�4���s&�M��0�پ������y��C�C������S�m��@(ɼm��Ӊ�rR������E�����h}�+�z�T��m����[H{��;���P������N?��_-�l�4!�e��t��>��q��U��ZGM���(qQ�V�H�`�_#)��!.M������x�[=|G��5�����uP? p���m�����v*}��a�L��"��w�>�� �C}�ɿ������DaKۥ�=r��t�W0���-{q��=^������kwᣟ�����������L��4�Ob/�6i����ml�Y|[}}aC(-A�Q�>3�9�&��OK��9�Xl^DNK�5�E����1;��k]&U堏_�ؽLt9�7�~��/uMp ��[�C%ȭd��]]���6Q9�~�����:'ЯAиD9��9S���� r�+yg��K�"����R��` ٛ�Y��`Λ�����o^�������3�s����V�>����|&�-�b[J��w�3�˗4���oj<�eDD���V��
���L0�T��'>=?�(%�YU55�2��YYY���$�9��b�rt��5�뺫ղ�(��C�ss��*ɼ�3��h�lC���[3N�e��m1Z�XR�����,m�Ķ�6�A��������8��˛�ƥ�>��$�`l�BB�8�⍥5�I��G9�Q6m�;]��Ћ'h��B���0�������ojg��K���y��n�0]V #�x�����<�j��l��A �=y�3�ѭ�Շ���ɷv�ߖ��hs���٤�����㪟�jl`���u���*;�=z�@���C���:g���FJ`����ŵ���8J����i1ql��-�פ���ؽP�?��m|��##�wԑ�	���������8^݊N�E�94���e1�58�7�G���o�y7j>IL��b��8���x'��g��!8Kz�[�����x4[�e|J� � 
fDO�D1Zp���^ ^��<���Я�?H�bv�1~_o���s�l�XiN�C8\h �\��!�k��hz�TL��v�㚆��X���1�ml�||��C��K+E�zi�*�	���t�>|�M�Љ�ؒ��b#�b[��qȸ�ԃ	R��#Y;?]�Ϭ���9���[�|S8�&_W>��S��o�wOހ��L�����ו��i뮦�l����DE�3��_V>K��Ƈ��e����%({su������t����(�r�2�����o�Zl��cFk��e�Fe2�Q����ݡ/���ޙ��6|�yi_��X�@J��6np� �1�!��0���w��J'�7?����FU�<�������;�����7oG�f&��'Q�n,�����܉��-�3�l#�,vv����32l���h�b�p��ٓʆZ54��e;��N�c���* t���YX��SD0@2w�U��"� �G�h�1 ]������\¸[��w����1�,���/�)�%�d��c��z
Y�J��͇�yK0���2v뭦h��
Z��la�%ȧ2����d�����@�lQ�ޕ}�Ճ��c�6�o?��\��]p$���\;�0��sj%f��gQ�䵵�]NM�ii+f���92��pdOw�Og&E��"BB±%n�.��Υ��Ƶ��~22z3�0���RԠk�@tSX�־�>1'E���/4j�e�I��D�)��w� �ƛ􍩫O�"_��1�ی�V"±��!ׯ�����z��£b|!�&�[�⯰P�o�'�v	�7Ϟ|o�̩��<?��v8����o�WA��c����&���a^���g��̦@��*�`�=R�~�Ƞ"��nC�������*|F^Z��D�B%�ϧ3�6��a��Sų�aq��PPRb�hw��]�������q/�Ȅ4���ޢ{�㰼*J ��77�/��+K��EKH�`��ԣ���>���_͇,����⢐\�$���̬:^P�|=�r�
���\�w:(<]Ōn����@���y��b7�;����L��2��t���䲶���-	��:���У���2������O�J^����ؘ��*�̳ܥ'�`=�r֓�M{U�ӟ$͐8�s�4�&��}��f�<�����	~���S�nA����qK, �g������ $�"�b.���3r�6��5�"Sh)�Q���x���&/�a�!͐�o�R�Mr����K��Z� 픬N���c���K�Ӆ�q���xC���g<"����̥�ޒ�[��S�9�s��,S�D�1>�2	}o¡� .�%G��{~9�r�n�3�hl���U�D�V�������E�$�-QC��H i�
?�4��4�Ӡ+K]�(ח�ڪ�'�崯Y�ig+��h��`���^�E�=sbUus�ȣ�:i�a�0�xv�ܞ$g�ɵ���fa��";{�:.Z{��9��4�Rє��Qe���%$�&\�;���~��^�s�o���8��&������Y���lL9�/y2�����!��
o�
n�����[��/�p�|���V��r}�ґ�Hʾ��hn�u���Wc׾��1�%}+9Z:r����⚠f����tvP�2yc� �k�'i��;f\�P�MZ�h��}��n�({o�A����vTK|�7]v���u�uB��u`���k}*ьP06AHLo`i� m�m�7��C�� ��3�2��Նy�^CfT�z���ң���wtFn��[��&���D,��4�'atfI1��u�QQ?a�_Z�I]$�n�%%$DBBZr		X�DJ@�KZbAJ�;�[Z���<�{�(�ߙ����\3�]W�E_�f��|���ȶD�\ ����n��]�n��Q�v��I���R���!��d������^8��cWQ��ǚ�2sxA����3�E�v��H�m�9+h
E�1i8m"�9v��		؞�Ab��;X��ڕ�CH���3�y�C� ӪB�c|<O����1���ߚ�c̴p�w�}Yo�JC�`j˙�c����1����y��L&�QaJϚ�p/��1���e�z���=}0��3'v�e��m/����R��ba��%��]���&��A��G%7��BE)\ ���ippmK��ԩW��#���ݨ�/w�w%(��}��$&z�Cu�d�{c�!E(�OZ�QK�(!&��a���c�<�oW9�$RTUk_6��̆�kTr�k)K^E+�?�9)����DT?E�*���vo|����R\�E�h̶wm�OZ� �D�Ҙ�;�r�D�!zC�	N��&�mrqޤq����[IK���Ӆv�|�&��As���p�
j�`��9��Հ�7��t�h��[���G�\R�9KMrJ?0찭(�0?���.��;�M ����;<��r&<��)����x�s��G�cy����{��N"�W�=�>CNL$O2c\"���Ӭw-�I:M�W�~�������H7��c���y=1�P���ƾ�g_��gT���d�>O�W�I�߱�O	X�9�� f���>��� �Uv�Pٚq���xWUc#��*���oݞ/_�v��������֯��J@�5�s���<��7o�r��EAFI AAHXX��tK��/�{��c�����'����N�>g{I��1e-�9��JKD]*C��<ٷw�Ҩ]?�|v�]&4��/�q)��%��F���D�Ndg_��Q�B(�͸v湔c��l�V �.,0�n�%�p��ؤO>SP�ǲ2�.��!��+e�� i(5777���ulfi9�~~P�}'����2L���M${�g����(��T.w�����
A�
�Y�v�_�N9���ۀ��۪�~m�"���Q�YO�S��8���k�q8��m<�zG�D�t{�2J&4��D����{���N�6�@ ds�}�B�ψ�♒��1!E{�>���P& ��)�2����Q���Ȯ�%+���4��r�6-�%�1��y?ŉ�2_�޲����h]�)/�X����8�n��(�7�	�wj��5�YJgfga���2�^߳�x@���R	�=��P^U�&�P��H	.]T��k�f����Ƨ`���'Kt�1�`�_�r�m^2d��ߋjW���Pr��w���o��nR�J��.�Z�0���l�F'�;i��Q�K�(�Z*��D���|,$j9􀗊�a�:WF��H�>&��QfJ�#I��H��F��咲�LN�	�4uC��K���%�3y���=c/���pv�5��Jv����@*0�����+�^�l����r�6�N�I���")Ca��/�&��l�p�;Gi�P�W�ء��ѧWZE��5�-l����V�?	�d�7:*�:��n�Z,}L'
`��~AшuRr�YQ�yΕ�$�4����aGk�x�Yb�<�6FsQ���L$��2US0��a���3�Ӕ]��;�|J���ҵ�11�6��ٞ�uU�:/?/���hD#t!��P鿻�[[v�Ҡ'z,��o��t�$V�u��j<�i5�hm�Í��}�ȧ��1�a�]�����C�E��S�����wp��ơ��.H��[yK�Bm_��@mc���mFA�G�ԣ���S��4.X��9��;\��/(e���k�|�~����$����m?�&������K++˷p߮�G����	X���߁����K'����^�Z�'���������%����&��h-�.��~��3�fŶ������E	�y��Ml�`YDI��0�"�I���=�c4��C ��Y��YrE�h�F����w���衪�ji�K
=HՈ���U���.Ԅ��E���Ⱥ-� �e���R�/[		:�~��b�A�h�}��y�Qe���e�Q�`�ޠA	jgJA� �6�3kM����p­��4E'R�&���������bP-OtD��z�̩q�V�\��17Q>�ΐ�_֔�]m�<򩴁�e����+�P��'>������A�U-c�goZ� L������ww}p�d`!�[f,}��G�"Zj���da=�e�K.�/VɅ
]��o545K��ZF��"�e��R��Jn��&|Z�$QkV2)�*�q
D m����DA�".����HH�Q_��5~���QC�u1�q�Ä�9�禦�Kt���U�P����v�gtyyZ�T�ޟ��百~�j�Pw�Au�9����R�`b�������S��L.��B4q[%!����[C�ެ�DV������a�� ������V��a�gZ�ӛ��wH�y{�����Eӷ���q�'Hě��C�-_�k���1z�T�3W
��!XwzS�eC��'Wwp�A�B���Ώ�ص,�媃��zlO>2I����U��W����H"��@Y�Pv�G.xsx� �&�e��qe����C��V��b��4�v2U��$6��fX�ǲ���G�j��S�}2FrF�������|�&��f�4�����]��$�{n���B$��b()�xDד�G�_&�5`�x�� MD0?�D�Pc]r������-�����±7�<���[Z3� �u����{=�����1�S3�,�E�N�"N"u��h�q�Jѡ�\8:x/�F�1>N~�2�T��Di��������d�O(8𿎅���!Q2����{;mÀ��'���-a��ꊞ̒��48�yg1�ț�B�G�}(Ѯ bMJ����Ev�Y�ŢuA$#��/����]����&eT�1x�ٷ�C��u���ͩ~2��sϹB<�윃�߄��������"�i����~�<<mX5�p���p1�N������St�!/��J�ҡ�y�B�ĵN������q��ׯ��ЛƀY(�gs%9茹���}���(�rI	[B�E��||��hA,V;��x����Ϧ�zy��I���5� �-��\Ӷ�A�_!��"d����<�HT+��I?%$�@����L7�@9�v�H-�8F�7+�0�
HJ�q"�Ǣ#r#���[�K�r��wα��[u���xR~��Y|�
��/��4^9;+�~�f+�U���ϒ���MX>�5������D��)�B�whg־gӿ��j����!�Z4���PoD  �.�%�.������㵷�P��9燤���倮��T����8������+�� �.���nynn����6x��*Lr��4���q�C��=��Ȕ�G�/$�+����pp��Eޣ�a�N�ϩ��ٸ*����~̐��"��=�it-�� [b�n�ǙP��es�3��A�[1���y�� ��n*�|I���\zx�=�7��sŊȧ�q�k�M/G�r�1AP��	p�؀��#�f��lC�|��&�g��cJ��kAI�Rܜam�k���t��+��췹��mx���y���H�����Ŭ	4����I+���ti����uw�^AUg�f�Ɔ�������*%���z���)&�<$y��;��a5Ů�i"`��6�p�۷�9&�߼y,8�}x���R����`�V�)@�{���q=�A�9����1~�Cf��3Kp?�lk�t���5���ݴt���ca��g�N��EK�D{�gr�4�Pw�A�L�)�M��D����7��5,>*d��9C$��� �\b�i9�P4��)�!???zgǝ��{Sn.9��#�����dƥvV����m��шU��	����v"���񼘥���T�V ��e�l>:q�X����������8;NU=�v����_z@8��H��B�
u<3C�!���)Sh��w���~�
�	����P5z�?�lY��~{�4�>�a'K��� e �ɩ)&g�啟Ɏ�s/�p�`1
�˷�9+H8:�T�����4���(̴�2�\��bm i]�{$a�GW��}p
��q����3D]�C�o�@�G�����H,�ǯ��sQ
kݱ�N������[�5��"�ìպE��[dq'|�A� ���N��-h�ꄾS�&��$;f{�O�����x��K<��:�~��	��"ɉ}_z�$�� d�@��L�R�����������@Xp�P�wꤪ"_� ��ީ��ʭ�ܡ���R����%)��u���� ��*�#w0��
m`P2 I�5�.d+./�sQ[�k(Zt�b'�m���f >&3�j��x���(��x�j��U��ü����0�qt��$A�ĹR�G �${�4WR}�Έ�gC-T?^����˺�p�|B;٨�vV��Le���>�z����Q�)��&v�����(�'�q�+�ٶ��߻ s��\)>	*�9���Ҿy
�#qO5�fgu�N/�@�2����h�JH��ZT2^!{fgi{�}p���!�pi���A� t���'��	��ǣ/�gR�@,���4Qמ��,7(����`	dc��W��x�,������6e��e$N/>��A�Y��g�B}���]N��
��;Ƹ�^�oǗ�?�[���\%Ʋ�O��y'��a*Ùm�FMNE�<������C��U�&�rƿ��T�(2PY�
�%�~��'�Y�5M={J'����'tx�Y�t~(���1�K��a���!M(�����ɿm�슺:�A�����yh	�h�J�}��E�@g�wS"��q2��1�~�������w�Vm��5:�<��wOMLA��:����}}�f����ڏ�1���QHzz_�`���)^%��-�}-�Gm{OcUa�<:�m~���ڿ-�_l���c�J�L�]�]���0��a�����͹��J�����_��y�?j�F3Kc���ҝ����=̿~���� �L���������ӽ���k��;���I0�f)9���=�P�B42�صG����u¡K�ّe%�,Mu}�u�\y�uC5 �����~D�mM�:`>�/��C2dga%'�h��C�h�T����H�5QL��Ԋ�3�,fh&�kFhH�Q�����|�`�JՔ"	aYB�!���e�NGO�(3�3��H��X���Ã����,�I/u(�H↕���L��;��Z<<W-@�u�o� #j>���q:َ�ۋ�s6�����ϙ�����{6u)�J�b��S/�<i�{"ԗ�2ד�gO�qN!3F�"�gͽ���H�A?�G���z������n�����X���7�f��;CI`��R$!&�}�#��5���,���|����ÿ}A��k��BܠB_K�]J�>���|�Ƅ��+�0����Ƣtܥc/��N���EO�HJJ"7p��=�&T7�0�� `V �Y���ȍ<�o��x������:ߠӜ����F�T�F֐u��Q�г���^
���B��+ߕ��~����6�����%��b�D�O��?<�:n��b_%�����,�da��4����A�2�?�D;�!�"�zN��l���w���e`����!��sX�ݺET�75eLYO]���j�ϩ��C�iF�r�y��Ą�ë*�� rRO�%�q��0���S�D�^^�G/�n�_�\"'�:��Ѻ�Ǒ�W�j��a�Z��c�_��r��Tw�74��چ���e 暰����E��0Gs󜃩���ة�Ci\��ӑ(�D)�q�Ũw�@�����=�;}�vƺ�/�#��LY=G�D;�G^w�տ��zT�2�E��^�Y=@�RlA�X�9m��Bv��mܴ6��^����G�΀�����zc;�_9�}�w�� R��Lsy3?�o���z���2��"����G���{�7�U��G��e�����GJ���7��˦�W�/O~��T<�������53�.�3�ݽ�?7�1�V;i`d�owo|2L�|�&ܮ�gX�5��aYM���]7������*-7� |���Mئ6�κ���Y�� ���������u;�a��n<�鹈0$����$��(#���yP,*&�ے�O$� �OD\\{Tm�VГ��!2&�n��f�)Υ8{e0�G���1��9���U�`]/���*4�Di��B��(=v_����DuX25�-�}~?�w.�*_�t�|���ҿ�^�dT�@[�4�â{#��bLp�0�#ͅ:F�6�2��v�,�@��t�w	�k�HS��_��*���v3�%���r���	fk{;!11���J�j2�e��a-)��<uH�����u�}��ʦY�L��Q>8rG�9�����go5ED��쐅"���So[W�܅$nm.��ٸ����4��w!3�Au�����.i����,:h�khK��z�� ��d��g�Tl���c�^����D������Z�.�A�7*���٩|aC����,3'�j	.��� ��O�SD��0�=E�^GS��=�G���eф�oOt��\��1�>����Ժ���6>>�/�)�x��o�S"���D�����q���G��_�����&&�n�F��NN���T����P�a���
���˓���j�C���J5�i]^F*i
�<֚�H��z+���<~t�\,d	~85�rU�[E�c�I#:�a\ҕ�^���w�S��"��n2���\�H_K.x����Ѯ�꘩uܿ�9x�9ã�1+��j��S|6o�ϲ�]N,��#�6������j5V�hooOQ����sk�TPޟ�rs�'��s���� Ǩ��&T[~t��[�w��[��;��N��4I&1���D�����TUUU�r�T���WL&���h�p2���^)�T����{~e���cCm���^��p�X��ؽc���Be}CP��Av,"U�Ґp�Q��'������j���6��C�Vv��d��f�Ys;�"���q��۹o|�ds�<�Tߥ���M�����6����\�y�9#6��u3�J_�i4�m՜٩�C�t�	\^C(�`z�l"RRq�D����;
���HC���%M�36rr�E%��� @����vya#�PZVF���3;��9�s��LU Cze����X�-l�v:������4�L�j��շj#�N�L�����k��2��X;Kxs0�m�]XmU�8������0�'� p����ё��津�/�f���yI{�qs�~�"���7"�ƾ�fe�t���w���s�@��8�8D�E����ͮ���!�-��$M=NHDt���٨fEM�����Tt��}��	�>'�XQ��N���2��@lni�`��M}p}�rE�g���h7;?��jJg�,2*Jy�1��T�z	�^ѝ� �Xni&S&h�*��^J��O ���J�&����\���r���#7��|Ȍ��w�����`��W�j������4ў���U.?��qV���f���r�O�3��^��g�F�����-�yo��E�j�2�|���Y�����뫢-�O�1G��0��xJ�4�]C�9�~^*�55š�q�4����!�8�\u�cz��N�s��@�pZ�� Z[Ǩp�Ow�1e@s�o��k���oY�-���0-7��ָeR䟷�O��lR��}���տ��j�#8a{|痥���z�21��������U	���/��X�D��"��1�� El��-\�B�����p[S1Z����:����M��DDj�%��p��(�*��X�_�tu)ߥ's��I��:���[2Sf\ƒ1@������Y������\�#@M//ԇg�^0f����9dM��xT_|�hf�9'����,�K�p�jX�ƀ�����h�5�tD p��V�ɟ�6ǲK}y�Z��튴P�=�\
�_�|����8N�ԌI�
Z	����}'P���O�p<����RDտ�l�s�_=�9��s�����ί�_��u'Ya��c�I�Kc�@��f�5�@�(��x0��@n(���E٢
�t�ڟ�Ϸ����-�m���PZ|�2f�^A���H�DH�\-�
}�T���o�){�sc�=�(S��mtV�@�YEAA�|�z��S�k�ȶPw!%֥��Ԗ?��^�F�X
�JH���
�!���rk�:�OL|�HR��ud���+2�y���Ge���&'��hL$��E�x��%ڊ�xE_� =�Ϸ��Iwpa��dnnn%��瑸8^b��be�8ii�QMǋ3#��h��xO^mb�����7�P�q"x�{!3���b��ͱc��2<Y���մ���ӻ��Z "����p��_� ž��-���}�֌,*��G��Qn����j#�u��ȕXy4�:�08��9�BL��#q7���)�@mt��zBh���89V��E�P�6�[�4g�kޡ����U�z�v\����%��j�7ul�ʇ�{�:NN�5K���_\x/��o7V�Q��#ub��Qb��e`�X_O*��ulfcs�q�i��ti�2�䕵���������d������3C�Q2yP�O����Ԃ[���s�٩;�*�0�G��������-�;dƜ��bn�d9 v�pg;���n��e�6R7�r}�'M�Z��"�VqIު�A|pi �X�ծ%dsj󌎮��c�TAO0��\��5��w��Y�n�$2���m��>\�-R9��s8U,�3�5x���lh�:�O��HJJ�E��Λ�N�MM5�Z�GA��J��r�m�}�������-,`��ᬭ��F�˝��.�ONO�TA�~��upV����-�y�a����=�+d�P c [�|�a��꺲�6��R�:C�$$����#��C	�� �OH޾v5���Y�Q��sE��ﯭ&�g���V(t������vS�0�(�f$ԌpPr.*+�~Ґ�s�����;9Ik�#E��~��
�S�"]�]ABd+��g�sk��)h����[��)J�aSS/l��5�fjˆ�(�����iiiI�u8_301=�D@c�He�������S�G�X���Y\�~J�Pg/��oQ�,ꖌ���u�R
��N[aDd&t^PAJUX6��(�� ��a-@>p�_{C���$�)�C� �����t��n��&�Ǻ�����	*���b���ʵ,�K�[Ā�lC^���=wuq!7.��Td�*�88�y)��f�����f�-l���!�n!�伀����o/�yh,-'��&dJ�������mG�T11�Q5G::���}�O2��!AXR�#06���	�O�x�H�_�EQ����Z�NVl�����]���u}C6��hQ�aD�tC�
ACk(KSk�-XN��P�X%8����ǖ��ƕ%D)d��ʶ
|�2�痒"�),`��E>n���&M6��y�!wWm����=T٨߽����(ё}�C��z����^��5��w,����F��^�
��s����j.
�J��D�٥�f�=&���!{���h�4�`��^���#V��.\��H�h��dB 2�V�'l)�i='���sm�� �5HK�4�@.oe`���m�o肧9��r�R��3�qK6�mŖL�;�����I�r�<˶Q�t���F�����*79HyUU���嘝��F�A�'��Wԥ��i�`9}kK�_E���$D3K��|gbb��$�;H�⑈"66��_�پ���"6ddd�}���� :7�)�	�diPto�+����<��2��;�J�
�Z�!����zC;5$/������~4�}��?�/KCK/��;_�u𔑬0��U����5���(�����{F@$u'5������#��86�sGl>��7����qz.X�W5�B�vxH�tA��à�Ya&i_���t�7���5�l6�yÓ�<�v�z�0ӆ���:���ۻ@��P/! @��8L./f�u;��ʂ��Φ)4���������mRfd���:p߭�^;<|�V�b������\��O���������� upʌuf�yVC��[�5
�#J��(ɍW>o���~!�<<�) Y�<���S{ֈ�����W'�2�P�K�w@ɺ������Gk��2..�YJ���Dj(�>!aw3P�&��^�.#L_Зڜ	"�����GrS�O,�D���H�J���x��-7��#�;7==�S����P���uC:��=Bxt.�%qɽRD@�{VzG�3���n�U�����0���?;���ǘ��PĴ�;�k�{"��_�=�P�걨,��<e�B��H*p�#��0�&7ϧ''c|���k)����И�w�����閉��-��H(ѝ��j�*O�9�l���sC}��Y>ŝ��2�P� ��Eo�X��,�w�Ar\	Ǩ��n�P��n�����#�{'�q�i
x�"�kw���Po9Ц�;w�p�C�h3�(��}����ZL۽="p��>�u��ֹt�Q���o�[X���=6�]���X�[vYC�usL��L#Ξ���<I�;A<�<�Ȋ��A.-�K�C���L��Ծ/r�1���lz_�����ϟ���>T��K�7z��qH|����"ןZ��JJ��U ��JHg��}V6�����֩{�S@m����{[�l�!�lP��PQ1sV�ꈀg�z��gB��Tb�a݈�n�����Qc��S(f��8���RH� ��%��G�zL4� ��篁� �J�<�;���좦�ݷ���]�Aev)�CC����</�����W���'''9(V����O,U�ʝ�"�W�ܖ((�Ѹ�:=gaa�?��:6��sZ�zX1ݝ�{��o����Q�YQ� ����Y�4�B-@�.���rP��OF��L�E{2��+�	B:�. ����2��6f��L��z=�>I��,I�~��=8a #�ũ,�}fu��Qir񰶾��ݻ����+.w�?��o���:��G��Ȉo'�.�a�d�%�T� ��T�`kKg\�+^����)E���ghXL�g"mȐhHw��7o����w��[��LMɖ�>${'���U"*�x�����K��9<:��)���m;+���(��)i��p�����(��M�f�>ًv�xs���H�!��`f�`F�E��\U��>�--v4obz,���w�I�����Ñc������p���{�(J�c��G���-}C�[\m�Z��f��H-�[I�"�gf�il�>V��uϰ�Bs�33X�RsS�!Ob����gi�N\\��c��b8:���ݔ=����͹5�6O-�8$���/�cьw/������<�KNa{X�-��8�s%h �Z���E*b�>�b-h�R�W�*�fd+�g�H���n���G���H��������|t��!��5L4�B���dRVT�W�KZ<��a1�4� Ղ��<��@R-��b��(�g�|��</�fo_̯������o�wx���7���Ŝ��}� {���K�ȧP�a�H���A������]02�
��˶�R� ~Ä���9.���F�d<�q�) ~�;�DJ>"t��lc�G�Y�o������1�@�
������?I�T		������{����mݷZi������f���	��p��
!!!�z(Ԇ�~~��o��G8J��4����q���D�%<����L*f�r�8������&�����v�5��iL�y��W�)�F^b@|����z�7HMҩ��W�Z;<�j�`�%~s]��{���Jc������.��c4BG�ȿE�k_*Xw�J2.6Is|�k�؋<�3-��̎.�]ў��v�����.>����ohBh�k�[Y�<%FtE��3��{�CJg��Ԃ���o��ǫ�+�؟�y�AtW �F����M|^ޙ��SS7��#��Ǿ��� v#3����Kߖ#���2��^&�%����^�2k�>!��`r�Y2����i�������[U$92X%�\�j
ME@���80�kWHX��W&��kݽ�¼��_ī�d��Ū��B"Y$Ϊ���d8��AE?�'�X��"�,�~��goo�4�#��),	�����M��}��<o��Ѕ�/i_��YL�����.3iQ��z6xǨ���?��-5ukx�d�XNN��'Hp>=l�ސvp �,xm���>(��e��f��d8�PYu���c�6�x�:R��y7}��±E ���������נ�5k�ڋ�ZE�p�=���Q�,��8���p���1U�YJ͌�L����w3�PbW�����k��«ޕ�\�h&����O�&�K����0b/t��o�QeiCYƮr��j��;��d���}�&��u��7�^�iq�o���,�)���_N������g�E_��W�b�$�I��ژ��m���&S��|I�uX��l���� \YˬB���]r�!7<�D��ǊL��(T�~��[��Ɛ�ɵ��(�&���S�J�nn����o��>�{�:-���U~{�ny�^������m�XTT���/��Sy4:���Ξi*�=,�^<�:/���'�H�������6��ϮAv;��?�0ߨ�.go�yV4V�|%��x����}q1��-A��@����bח��ß��,h�J����뇷���kƏ�a8@��2H~�(U蓪[�-0�=�H��!�������Œj�-52��Q�`��[��Xpz��F��v�6Y�
�6�ф��,[O�g���i��B%^����-�N��wBd����X��y�<�wW�� {V��nDV麘m�q�5nM�Ϧ-Z�$����s�<⑨V�6O�%9jr&P�&ED�7.�VWq�"��G�gml�@m���ojo����b�:�FB����ԁ>{��'����o�*�(m�K4!�q���d�+ό��>�7�~��9f�^Y�P�?g1`�Xg�% ���߲5TL�-s�9�E*��rx�Z�LTJ��7���%:ߙ��%J�}y�`q��u�kSS2&�|?�l������
J�ͽӥ��5�z
`���`�:6>5, Zξ<���PN"��(�g��Y╹6ä�C����&P�\�&�,�'&&-��#3;�
�G�rF8^_�O�V����^��=�X֥k�dC5|@5��g�EPU`�~�p����6�~���D��m-����F����j	/�DK�Y�kd�l��QV�gy��T�*w����Y�~-g��Li'(�E��U�Ը6<�ss���������U�w�
/dM٫�5�M+�/�?z�.�t������3j �]E����^�N[���d���!��\�.������&�+22��a�V��"־o��'>�a��D�<`M���cA�&?�I�-���jH�Iy��A1��0��,)��mSH��J�/���<b��Ukb�(<���~��̷�w�xw���`9:l���1hWFmʡs:05���׵e6tlll�&R�D ��[�H�Dr���V���F�����ӄ�.���Mhg��PR��?L�e#���Pj����{�j�e-�b��V�������3��1��'�
9���=���\����A��[PDw�4�$���ݼu~��i��my>��͙1�~),/SoH�.h���tf��� S�
��s���b�(יl4��$%T�Ы9�Ǹ�@���G�x`fַ�C:��Wmk�½4����S��|�K��/g������!�X6s����L�
C���Iy��naӢu�	���p����ŰB�~n��PH��dU�g�5&[����?�2jy����6V� �_S�9�&��&Jt�v��Hb���C�f����V�C�>j����p��"��/҅sD�޻kY'�19LH)_�}������bJ;\�]"g���-��j�]���!KYYni���]d*n���c�(�w�����-˿}���nm��K��E ���Rq�y���}j*=��{}P��] ����Ĳ��û�s<6Nf����[��E��-Ȟ�e����R&�H�%�}���>̀ ���c�N�޻���[Yy�ߦF"�@$���1^Q���wf{l��zy�Z�	�N��2cj�~�%�r��Llu..~Cذa��=@�:CE�M���ٸuJ���[y�!�`��+�|^NN����aY��Þ�cçD-�V��w�� �}(렙@Y����Z�ų����u�v"��u��->�gu���
dj?�ɉ����r��9ƞ���~���[T$���zà�(��S_��tsy�n�7D��q����o9�����T�>����Pr@���X1ȆN�E��0���M�PyJ���_��p������/�ܭ�P����IrR/c;��09$c*�&��w���)�Ԗ�('%>ж������{�������\��:F��[�r7�$�P��o�/���O��9 W\̝2�y�U�Q;�x�j�nP:J�IH,�`��/T=^�wp��uμJt�D��
�������{<R-$j��*�*����,�*b��N�B�������HYh3z ֐��)�ƵϤ h5�����A��Ik�Q����e0�3���(�""8$�I���1�����I���O&������s��힟/="
���}�����d��'��&��2�3G�f�0����s;�ԉ�"
2�4�ƀ���Tt�K0����1S�1qҍ�=��r�Łv)���O>����&��66V���C�e�nP7gޕb^�	�'���J���IDF�fs83ֿ�x�&�7d�W���~3Y᧞�=��n�('}S�f�h�	7<�Ƭۈ��H�P�gx�c�Y}_�j֜]�(����cA2"pp}%��͔12����
ä���d{q����HT"]*���[N���w@r����1st���[���NJ��㶵���w�(�O�A�:?��U6N� ��|Tc�S zǈ�|�J�!Y�zidA�[9����.�:��i����C���!a� ��b���^���=k�nQ{������J�s
Yḵ����8Vm93�P��{���"�s�wN]���)I����������6I�x������*�r)���&���ܜQ�����ty�j�`m�#����9��/}��NO�+�]��/q��7,/��v!�v?��Ս�%���vpP�����\@�x/
�Q쳖�z��*�Ez�* ��YX�F�d�ۀg�E#-,0<,�030w����a�,!�}\I�4ᵶz�Ū�`�Vʉ������bh$�О�
�_Y�42������+�q&�i(����_Mv�9(�F����mU��}Ͱ���ۃ�G���V(m�ti��� P��!h\�:IojlD:]0~!E���:n�N�a�����I������8�z�A���>��#�������c�%ķ�����_�m]�}����p�;!�f�#S�u`:f	�����$�Ps'������د��F~b�a|�-��Qm5[j)/�p㖿�Hc4`Y3�1���F�iio6d�~����M!��l�-��s�}9���c3́%Aei�Q������5Z�a�ݯ�㥩*���S��SSߪB���24�G�r_�[jk���I�dƠ��"2��1���{���n�'��|�Y�MSG��jo==6@J���Sc�M��7f:���MG)�B�v��a�Z�K���׺�z�q)X�`�`�1�-[6��o���=�Z�+ s3Z\�rKOO�_2eF_Ǿ�;��G���O�.�"��Ǌ�a�,�s���*[ ;��j���|��4uv���D���4�q01$�O��xđ0+oi�r�%�|vky�b�����sZ�:����}����KY^lH|�6��&&��`�FCTl,��g�����YC���zC]�$�y�Q���l�����-��H�u���`U�����+�����o�4"��6@�������k@��$M�}.�����]=�z���𜵵G�=�R��2��Q��B��[ e_XJ�bAcctoo5`qqE璌�"�����G�u�<O����HP��d�.���g�mlp�rßqS.�_qy��p��l��ݻw��-
u�k蘍��oP����۰�����L���I���F��� ��1������CX9�~�xP6�B9tSJ��i��rI&�l�6Ǣ��>�4>��O@MQ�AsRs�u���8�8�s3O�
�{�=������Z����w�� [�ҴGɮb���t8��_�<���C�����~�nm�e���z���Xq��@[�A�'50@4`ř��ϳ}���%���C����v�]�2,H�mo;y5r�남��9�ԝ��sQ��iV��'#�R�"�*����.��X��i-�AFjI?�z�o�ߙ����
l�J
w���5c�e��>�7��n B�Ʋ*Ԑ��U�{�J��/��{����BB��Ռl�%i�*�)zn���}�
�~]���ORj��(՜.Ob�L��}�^�]JpggHRJ�.��5�B;*���6"��p���9������U^���S�r��(��	4�"I��k�q�!q����bs~Y����)�B�6�xꀥ��C�u}`Q�'�m�0;�-� 8��]&�[�S��P�x�nR�{��:�� d�Ø���)n�ܸrK�0�o���ss�6s����;�s����C��h�W��0Y�QbvvQ��ႉ��k)iiHd���=�&}_?AB,;�"��8|�l�[ظ|��J D���|������-���9#uG��ffO^h5�;(
5��^�W�����Ĥ�P�N�k۳j5Rp���z?����;�� �6P.�s���5�-��8e�}����xJ?�ǁB��#�6�g\�q�!"b?+ ������S��x@����%/}n�M}a�9<��9���`�6���~X"3�iJ<�|D���������I��	K���읚𑍎���j�sߵ8�]]�Rɭ���X�]\\|���a ���$�넪��S��z��/(�jY��|��C�`s�����&؛E�����=A�D�*��}�"���ރf�v��%�:|����Q��QQ>��0 %��t��Hw�,��! )Hwww����,�%%�������+ҝ>s��s~���⸰3s�ꚙ���*��8�&�y��{�y��s\\O�6�������1����j�����e����0�x}�����*I�۞uNd�ሇ�w��W]�[���E�|�+Ra��G�iL����-�.S�1���:��8��+��:��������K�3����"/���+��}���^qo�~|��X�}NsɝڵYՈMz�mN�K�m�����tW�B���@H�c%��"n߾psY�qޙ�$GF��C���`��]n�wv���7@��
��Z�7jǿ�Dx���ׯoQO�-��[��� �R
�����1�p'L����ZZX��O/��r��5= �J|!�7�팋��+��_�� >~=�K�K]O�ymȞ�Z=��E~I��e���Q�7��ygg�s�7�888�E�q��u��}9��_��dC@D��*-M�<��0� X&�zC��jO�e�80��i2�����H�߮�#Uw)2�{b91V�c	��^ ՟rQ��*������Η_HT�Z�6�;��ݝӼo�;�v����o^w����PQ9a����(
�}wP1�T&�
+*j9n:,2� �RsfR|�
�W�O~��3鼕<�`i���`���KY���Ip����c��������Ze�����I/�V�z��WdB<�,�6��(̛�b�w
�����cE�	��1AЇ����:le�p�����TRq����F��跉ec�;�F�1��������o�b���Љ��m�f�D���Y�����ֹA��(����yN�|�53q�e>�͈�s:��iЋ�x�'������	WW������A���G�D�L`#Ƹ�(t�@x��S"�uV�+�����1��H��j�&�@F)Ϟ]��*�B�I�%;O=�H� �c�H�Nc3�|?x#>�75����	+�
�d!|�ǂ�����?���;R��r�E����,��g9x�hV~��002����5R�lU���2�C������� �C�:��ŷ�[�t��I�С"�\n>�`d����@Nl\��~=0��������70z���	�ۓڕ�/���mm��{Pcٿ�����&��\Rbj������6��G�b�� X;����m^dވ�y�ų%Z��cu#�d��x��v�M��������^���m�s���d�kJH��3Ux&��,{�~�=�����rdك�痡�@[�T@ۛ�.;j��9������趋}@��q���WH���ncj���t���"��vh-+k���-e*#��а�����?�XY|
�h�t~�� 
�"�����l�b1��"Ɨ6���f��m��%�\�U�ŵ�4HY��������u�5�t6a+��o�j��b�;����ȝB�X����'< C^��N�§������p�^����w������W��7	
B�t�<��w�~��_G����̜ǭrh.d������$b�#(�:��ũ�3������!�����:T�(rپzl�����؈T�U�MF���`GEv�����冷iS�s>z<ݥ���v�×�6����=Iu��do��K����h��P��y���hu�`0o*�kn"Z��Ǚ/���	������'ѹ�|v�wT[,�*%���5�"� ry
��>�(3 '&2m]]��p�vMLp�D6n}�R��k+zя=��r��xe"?-5u7`�����mͣE4j-����6�ijn��E�^	�U(��96�NL.`.Ҹs*!�c>ξ_�@H�-ͿΥ�rs������%555�D���k�{���]w�=�i��B�0FX�>D���f��hb�ͅzyLR�l�=���Y��p�'ė���Η�|�Cߵ��>�����Ed�ںF���Y�{Δ�,3�)����#�wAM����Z�Р���^��ii�z��������mA�I�I?���}��n�~F;�8�ba!�/���{�ϯ��x��v_�+�nb9��GD/�w�,~i��X;8(�N�hTUW{�����&�x�����|YȽ�w~?AP�%r�rE����б%�"1�ھ|���] *�1kZgD���~,OE�0�}�l��C�g����~V���=���&��N��hK�LhK�5�<��.u:��KD�HS��)�"��oW]�����4;�dI�|�R7U���z�֔�:$��dm���ǏX+��f�<��~���ܒ�e@ 9y���
 C�X�������_����� 4�y��dNd���u����{�۔���s?�-�A�����Ò��yv���������v���cz��O��fr���f����^K��k���)��2������$���p�Õ��4�IW^���W�	&	��7��g6$��­���]'��m*3${���//C斗�Bca�����>����Eo�l�P�|q�ւ5���:J, D�R��w]�u����ggPg�чJm��������8���)�ôFl$$��ղ�ˡ�Q"uMM�elXᅅ,�ĉ��}+}�C-�HA�qS��qHk���Ņev�� Y�3�bVNL��⼕Y�3+|�?��~52ӫȷ�{k�L��lJ���8Ą������_=I�x����0a[��.U�{3������\���-����PfH�H@SK���f|O�Fsy�h�FUMG��v�(������w2�|Y�!}�O<=�
�KQ����@꣓f�&"&~jn��Ǝ+MEU��w�d�$edꌴ��avT��@g��߀o(*%�|y 2F'FKCV������IDH�Ch�+�=����𹶨g�b���.Y��3��}��q�?M��|�u[�y>Ҋ����N��<�(���	����e�������,@4�
X��	
�:���ǣ"g�[������K�����XU�0Hs�'����x�,oim=�w۬s!�����'�/?� ���_��.��1��%�y�%)yiy_�e��aY5'������a+��:w�Wll,do�9Ҳbt�>�R� /���G�����/��L��$JJ˼���A�gV׮-�=��-��^�.����~�&�� k��K����7�r2q',���[F�'8&~�_V��[^�C�dk �|���e�Lg1���;�Gw)��v��"��9���==#��nWyHп�I��f?6����H*����)_&�������#��O��?AY�:���+~֘�vD�݊��O(�����)CCFĦ�'q�	�ܻ뉰\M�9o}����.�������)I��x\�n���];�(j#����U�R����Q,狭d���ֳ�������s�C���;��v˥F��8Cq���	:���DuWv��;ᨯM*0o/C⡧w��?��Ȅ�T]�U�	l�z��%��'���\\\���%UkDe�{��&�0ɩm @�#�ĩ�<JK>궎��i���S_��s���S�hδ��1�F��2+���dm��PVc�t�l^>���<	��C�È՛j����ن?*�����{p�-�9=�Gؚ�v��e��++lm��G"�YUĞ�Ƈ�6?�
u=:$a��
#�ĭV8�B�ry�C)$0�龮���`�����V;k}�o̪�����w9�R������lh�i 2i�ث{��*F�/.f��� S�P�
�w�y�V��b�[��������H4���.�y�H/$�3}+���k�30].����Ε�����נ]����{����z�8X����l`���tTҜ���3�b����%?���@��f)Xb����? �#���yh֪s����$��=э�[��~�`	dO����q���'�d1���Q"�=/�~����d�a���uT>�1��	 �9������:�Ur��;qp|l��	��--�^�f#�����[�hSp!˄�7�'�.|��hl:"X��fb��P���Z��&Gk����(�� Sf���
��-���g��d�!!1��1!~�����R��u�W��֞��1S�얠�t�M���d��M�Y�p$��Ry�#�"��j6�P;wF;"N�Q�&���`��.楫&�遊�m�#'#�9IB��fǖ��[��#�/!��QmR�=_�ɕ8<��R2��M%�Ð�lEmdf��n�9��#� �%L�/�!�ZŠ�7���e���$�Q��a��ddf�%  �������{����=_�I���I�x/�����8��3o�æL,6����+���
1YY��v��<y�����.��u�g�=v/���KXh('�ꪛ�fm������W{�#�mZ��阙'N ^�^0���o+�>A�p�q�/�62�Xh���WM��R;��:ڶ�Y�n����NM��@����Tѭג�,�~��Ti�}!z�`p}{-���9Osi��Xz�?Yii�{wщ��0S>�&5�D�ļ�"��?P�W�8ݥV�r�g=?<<4>��ZBp"�G�B(`d� $q�_9�@|z�I�v]�E�ynz�I����؜���ٜ�+��k�}
�!���Ǚ�0/0����m��6����`%���qP� #�B���4��� �0�<�	Bb�=�©��o���Q�0-�4�����>��7��M�ŉ/;����1���mϬ ��WI���o2>�q�K��ɪD[�o��������d}����݌�JLL,i�@���'޵}�#�Y�������������zK|覫�����Eж��d'|%���)&\���dA�U�'�83a	;r5��Iʇ��Ȑ��1���lП*��rH�橵+�xP�bc���-��ٯ_�y����wŷ���>7�61<���h=�J�������� �dȨ�ػ�3���?� �>��Y�~�CL/�a�$N�|�i7V���GE��SS�����#�ohj�C��Q2cA��J\�Ѯ��']Y���w"��L��eX��=*E����/��*%��͝�����˗���|����-,��#����^1�mE�>�"��@|Q{h���#@�>h���.)-+�7��|����0o4bO�y__��49S�t�&(����
2'������QT}�� G�_���eI�������J��o��۫���.1>\nmͰ��mE;���;=]���!}�)�1{vХ2�k��~���pC�����O�:�}_On��V�'H@Q�jAs��9t��B��Ԉ�O���_���������"��>^��a��_����e��z�
oi�v�R�rM�VM0��*�kYOwoo��svZ��:����9A����#g��r�VV�,�?�Rc�Gs&(��`T��?��J�Лiq��tO��}�����Vi�y͆m��-t��Z��PR2v�z^��k?{F|��DDB� N���+�� =}���7�,����o�Y��Mo�R�~_��_׻�~��8�`�!/�z����OS���2��<5�3��8��z�$�ܰR��9{i��Ü�2�a�gK����d�6��Z�Q�Q�UGp+�#$Kޞ�.�e�Ff!Q�zr�A�����j����1/��S��ՕQ+_&fv��NXNe�8��$u����#�Y�P5���^����>�<Ɂ.n4sQ�,1�rRXC��:�cbrA���^�Cvp`��;9_&��9P�}��;y�Ԅ/���,�#5�w?8<���p����%���~]ږ�_?�h�IB�`b��e��i5=�'�
O��k6rݫ��翺��5ƌ�49?�｜<��^$"���$�Ǐ_]�Al~w��Z��-B�1|� G>��>�&\����^�'�6h������Z_�*o�/#�7�����0VU�D ��O���,��S|d�ӗ�-��w�EA �PRQy���l���+���Z�ww=�[%2�G`��@���$�#�͆��{�1f�jv����σ� f���l��	��8h~�������W���5`他B��I��O��i�����!����=��L���(��v�Ŕ�/ŃMe�_�.	�JW_����:.ٔ�
�wk���׊�S�JEEȇ���u�u?��ؑ��.�{�K�/��"�&!'�;z�X:e9�j�����
��+<�IAaa�*������i11�*I�a/��-�ϭ��;��t�ﭜ���t��j�s*WCg��*C��x��X���Fv�����XV�16��[o�_]�4��Q���Ȓ:����_o�q���-�utxx�EL�y��[ޡ��۶���ᘥ�/ֽnv���P�w����5������^��2w:��H�4����(zt��A*#����iq�>yW��n���%���/!�����P��v��3_���jW�S�|k{RGmʷ���OA�tR���d�UU�� O�Y��_�nRi�?$b��ikߌ'��g�V��辽L��MD�O��N��qS9����U�[���k�f�پi.��y��<3�Wq&O��\ڷBo�UL���[<8B'��s��-Б#o��X<̶n�t;˻����FG
0z*��k���X8ן�����0a���Ne�iAp���i�g�k�uz?�\�D����z���Ȓ;s�X~������h)������[N7�	!�2�3��ٔG��u�K��+5��۴_"�����|q��'Yn#cq��h���9�&�<��۶,�r�_��`Z�c��e}��~oo{�o]c�g��Ǥ�'�09�-��_�XA����;��q�����C�����.C������#�i�_�n$§h	q�x��N�Y�C��ε�U
�5�-&�C��o%fd��+���95t�,���C��NEm/�>���}��ݺӆㇶ	�`Fj�ɺ��8�Z;Z:|캖�,��܁U���T�Z:�K�1tOmO�GJ�^ּ�v�6ō,��5:\�g7�;�T�/�e�++��]`t)*SssV�k��X�}���Ԅ;��	�4�T^^^Ō���II^�*��-c��"@��ו�M��,0d�3���42d)T��vy��F��)?��S.8���8�v�iX
�|u�m�ǚ�ƭ��C�*�-πmQ���p=�u���}��N�}���l�X�߿��<��yI���Q`������pcjB\�㭠�B�I�+�Ծ(���ۆ�&����ɐ�}�'㵡Q�����SW�%/��;����umE��m��^8�8Lͅ��(q�mk����N�.��4���ɉ���Ӗ��[�LII�۷�i
�x�^�gO�L�M�;���7]$�w{%�GPay�v�S���F���I02��@O�.�X�Q�#E�[m���r��\OuUA�����Ɗ��������4ˁ�U*/���bk=�]�sPz6��io/Q�:���R����8;�#"Y�_�6T'W�E�?$Ŷzpr4��p��ZTzv����un��G�v�򜁞!$�$�"st����3�4)b�#��XI>��&�����=�dqi���������P�{(Ԉ���Ü�5%fR��~��$Ԧڋ���{,$9�s⯢'7V��aK�_ZKfƟ�9ã,LpP�Z��\��Ɯ����&/ػ����B��OW��n�UVpwK�&�a�ݽ{7�R��%Tij�ǃL��1�Lx��+MIONL�&��|I�-�v^n۾�:��Q,'z:ha��2K�S_(�sm�%]4b��Ҵ�����\�@�s!us3�������J�&� ��ޖBG{K9k}��VAߊ��x2�8���>�S��!1��XS>'�}+W���\;�
ޏm5d�{���(z�1�9� 
���@�<gG��e�9��L�8�%��$��#�k5ߓ+6�aJ�[:<���		z�& +Re�� {�W虘4H�X:9��L�{��RUe�y��-�Ք�����\��d�,��l6wv�����H8f'���wp꒻@��Pe��@YdH��)M����|�(��J<
���(�0�ş���*LJV��jr�uVzw L[��o���
(�Qm�m⢃���l�]�e�ӝ(��n>p<4�ʻ���N��C8r}j�>�Aqn���a��g�՛�@�� ���%w���pVn����1������n利�?M���+�sU�PF�9�df�M)4��S�J���ȽŴ%6d� >�y���y�V#C8�.�%`�ݥ�&vf��ꠧ�LFkA;q��������MϠ1�n����3l+�\��-!yj�cx`�ɒt$�����DCs�� ������
ۼ�VRߊ`�Vn~�J)�=��z �''|��P��'�zm.���އ�'r	�$�k��/Eғ�i��|��Ԛ5@M�s��Y�i��=[lZ����(�_���㝜�N���i�Q��^c9�8�>X�9Ig�j�uQ4yP�$
j�ZX������z�$�yz��p<�o7�X�����+��kE����Bs��S����\+o��#�Ѕ������gdİ������軷� G$��Vu��x���d3���4�6%&����B��oL��$B��!��R�:az� L`�l�q�L�8��gr|�a"����B�	}����or���Ń�^��E%Q>UJ�2gء�]+9�C�����!���OdI��^��������B�q�x~�S�����]g���9W��W�Č3 vAdr�9�~�(CX2 ��[�x��9��0_`�:�J(mT�Alָ���xr?�gkce�)W���Q���n��Ut��ɟ-���$���p�Z�_C�w ~-8{���ϥ8W��7�(�Zh]�5h��s��u�6L�����ʍo�6���^QR�ԭ�����W�r��L���$ʏ)*")�|���911T:�v��n>mǈ!AO�1`��oN������H$^ٯ�DLJJʝ��L����X9�`*���-.�[�q���a��`�m��i�
�c�?�*����/��D����6�ʰ���qF]]��#�W�|t$�oФؘw�Vr�HijI���v�{K��O9h�����6�&K�k��o_�npa�d�I4��j.���y�)�AoR]�Ph�݃^BيY�g�������=�S^.���&.���(S��{�u�l�w޵�E}z�F��ٲ�k�N텳�����Z�w7��,�7��$Y\$nT%�3�����	rG��wg:ն�����ǹ���5^R�2`T���ٿ˹�Gq�.\d�W/������,��Y'	����(�����|��f#���($�+z��I'���=c��|����s0��	nE����1�C� t��ȓ����r%�@���E��qKܜLK\���C�y**a�����U��/nmz�>,�Cz���k���Y[_�w�x� ����15qJ���5 ]7���O��.�껺bT)B��Nl.Ϻ�E�HYY�t(���;/Vk�c]�K�3�.��:��M�[,(�?��p���[h�9�HT)22���e``�r݆��?��+>wp� z}X����iq�^}ش��h^� �×� )�j��s���X�X���"�]74r����m�T�=X"���ź�O�����m�g�������C,x�k�\��$����Ms�h�ۂ���t��ܰ�[c�PL9<�65?ˌpL��b��o�	#╿�ʹ�a��E?;��)�,;Ҟ����2 `���#t	6�XUB�r�|���e�v�h���JQ���Z/��+��
A2J�����,�{� A�!_k�աuw����T�C�_b**�^I�$�����m��a��E}�D��ׇ�R��8P��pvu���C�5`�4P"y�'�+��A2�?<%�iI����Y��Q'h^�7�<��gfEX����C8׽�2}>ޡ��ʑj�Z'�ӑ�]��v!
m��f��^V9�����F��M_��{/���� R�lRbE0�\���R��^$ҵy��N��67���罽��L
��ϻ������뻏�b��W��B��N�sv>�z��-�5��vQ��ܹz�C�׮��"黦&�)wz��%��Y�@�)렐��8�
�>A�LgX�$~���~�s�}ޤ�ö�~���/o��U�s�r����T�#֒�l�JTc�	�����'�*��k�J|.����G����Ax~I�n�m�׽��u���OU��@���3���t��u]�G�<ԝu�Ŗ�{�;b�p)ǭ���ۢ�Ti:3���� �����]r��+���xxT�C�s4�Ss$�K(�8A�ڳgĜ3{0T��S�v���))�KF����N;<In/� �9h�(~��ߠ%FdA�\'GM(g��|/0��	�Y�5�7�f����n�����Y�)eQ�.����+ƪ7\�ZZpl��We�a�)���� ri��|!���h���/�����T&y�v�z!�O���&ݟ`������32�U_�Sg�;�cc�X�I��x���P��E�����mY��$������3*�5���`��J<��T�W�� G�Ǳ�h�_�n;!ȌYҍ���tTJ���D׎t�UNn4��ކ߭��
���ӹ�y��;������o�h����ᑥ����P�B*;�(�����n\o%֡ #|V`��t�=rӗw�9�i�V$8�yT'�YJ>�יN3
��&���\z���؍���\�5��X�Y���V��(�܈���̥%�q�">6iO�EjkZxE�}�q�L��P�ߢC�5M ��L���-s�	��<M��4cJ���˧�T�=?=�ssݵW�n�ߜ���E��n�<���[�k0��a���^�4+P\��jhz�Ʊ)��R5vG��PϽ�s|T��[�����vy�Q�Y����;�+~�)Cs&��7�g?/q���N�O6l�<�̚�3hmmc�s`�Ά���X� �L�S�G&œ��o�ί}Y��I.������\p��"����ܦ�
.�vh2��`��=�$�D��}͠rV��B���� G�HD�ƞl^�7��
Z���������@�v��'u_6~If���u�M���Ǔ0�=�dk�?AFGd��qm��������"�ڥ�5r ��ÛLهa�**$d�C��V4,_>�]��p�=��-��lNY(+�-	�֝���6f|6e�����;G�|�{��٧���?�~�ntӷH���ō�l��O�,���)u���M&�%ni��$#$ͳ�b*O�[9^����v3!�B�:~�g^d0B�~���ntX'p%�MJֹ��W$z�$�w.��l���$��� ��@��I�Xr��u�L����i�����X櫻D��.�\�Y<`�Bt������.v/����Y
w+�J�}��jK��X��������hv��E}%��2�|*l���Y�1��ϯ]nj���b�u!�ܑ�ud����:1L�����.w[@ظQ��&��#E6���������3z���=� %�i3C�%f�x\n���b n?�/s0�����~��#k�C�+͋Py ��M�X5ĳt)�/����.��g,y�h�5�/�TV����9J�~-���J%
o`�ja�H��J��2��%߷�ɒ���>��o�����*ྥ�s7���)���c?��h)�,ʺ),1�f�3i@NS���o��-�/n��*���}dJ�F&ff�P�&���F��4���z]�Xk������g����v�q�l��߿k��;�%�^�q��CvlR���B��O��*&���UZ+����ţ��Q�j�2��2�u���@�3����Vp��Yy�"�`��}�]���)V7�ѻx��\�]����7�Z��*�P�X{x�0��]�I�W�B��W��-��CMY
(�_��茸W�a��� �0��ܵqȒ���m(�v���F���d��<^9	��9��Q�8�v���RҤ�wM����b�����㋶�Q���;�7�}
���=Ʋ��y�j��������4�A���{` ��\�����x4p���hϖ�'u�V�0--�,��»öךLƹ`�"�����y�:]QP~�V�P����p�l�X��l�a�=�*y�C��>um��Ζ�C7.��m)��7
T�N8�cI�9�n�_i@�!s����\�k��m.
��Xx2�@�k�I��U�O+�ٽ��X�cmӕ��5��o}s�og��Fw����R�C��#u��*�[�������C�]���B�#��֓�%��RN�^Z��я���Ε��x��qNw����>��UW�|0�=)�/xc�ơZ���ܵ�b6��\'h3��I�k�!$�����V^��~��
c�������j��Q>��M�И����cn"���a�Rd��✌B��
��Up�jR}��E%��Q%��ݠY���h򾿌霬R��p��}
e�0
����Q�L���%(���^{�_(�$ƈO���r���7 �g��`g� ���;��l��	�z���><�߂-Mm�D�և�NIyyħOr�s_)<��qQ>~��C��s��K��Ӌ���˼���au\w�$��� D�vs���8g����b{�D�!x߁�z��q�u���sr|>c�|���0�2 ��ԕ3V��:�ȿ������D�,�I+�n��Y��q�bہ�9>�;w�|_�7}��J�4����Uw	���(������R)JQ&_ �K�D�&ZN������2��h�P|\���	����g�2�� �����|
��_a1�͋�9�cu~���Ô���tR�=� �ߺ#�2��;҂2R���ߧ�V���f<�r>q� ���"� O��ռ=���lg	c�u^e���x��q����K�(E��XAPh�mw��o^G���.��\ܫw�fܳ�1x��G���������lpmN�"ҡ��U{af�������/��4�*^��q��K� _����5/�w@� ���`E` ���f���z �/3 -��4RB�����'論��7����v�Ɗi0f�uD|�{#����L�R��S����~on��x����2''����3�X�"'�dnb�=Z�u���\Hjh���ၗP!%%%�u�8���<����rU�4Zn�y�2WT�������P�����1'�Bnw��U�/�P��]���wA��|����:K�w��YYo ��6��/��mKY3.x

�\F�w���>��K����v�s+$m6�WR�l�A����ÈF����EP�(g�ZSdʷ��,~��3Ǧ'��F\����B@�?��<� HJ��F�돕]R8����&RL��Ǐ��4���USP�M���� �
=���F(&%����Ħo]þ�g�==��T�%��G{J�O͇>5�/ېZy:�0��[�n�ZZE���6qxH���r>�����"�g�6$��ʒ#+.�Ύ.p�>"��
Q���N��xk�}�f|;��(�d�����f|m�[`�3�?��%�GքMu~{�  
P�'��Ts�7.Ed���{�#�hZ��L�X�Dd>P)�E(`��#�H�gc��|���)��3�_��	��Wt�Zt�q\�I�bt�m����W�57���)l�U*�ck���d�!�zR["(�?���t��Y���7"9���~10��A���6�ε�ol���u��.Ri��+��_ �r����E�6�K⦣��ra�z����:*�wӍ�	Pŏ����:��;g�{����qH�t��\k,�_��q��a����'C�I�ꔷ�����ɖ�����#���s59I�x�r���c&��c�ǒa�'����L��	�vG�5w	f���[�X��?���@��X	�c�'�N���5�c_һ�̿]P�:��Ԅ�(�`o�u���1���A�M���d�˰ 
C�6egu�1		Hbے�vd®��� m�mw�y��1��JA��ً|��U��;���g��je+7���Fʙ�)�9>���(�u
egWW������?<�o4��t`�3Ԫ
Ş	�m�G>������z����B���ҭ<�a:��c�{0l���'V,rG>�黑w��0Nɿ�V����sJ[�Pr˻�6ƌt+�R�Ԅ����Bw7}o�e�z��[`R �m���M��e{�0	#x.r�^���*�O�O�d60���XPrz�"��J��X?��j���¨�������܂��0��@�֯.�`�P��ɚ�Yɖ˺���� z�,���#̑��Y�4��թQ��T�E��Ǐ?|ot�\�^Y)���U�շ~��8v�/��*�?��*EH��_�SJ����p.\�� W����z�5�N���fM�B��TOȅy�����*^{X�0�*>�+\!w4 )u�.���2d�J��IkY��8]��[��a����9������:_"+V�Z��/��O^/~���F&&�?���S�rk�*��L���VMa2 ���l���W���{�Ϻ|:B�c� ��F��EG��܈ݭ��?Fڋ�RC\l������3[2�OL|4u`1<�uj�e�/N��w(�E��Ӧ<�q��`Gw����͔�3�]r�I-���F���-�j�E:�IH��7.�82E]��_��V�"��*��]�9��qǞ�C�}@�tTY��Wj��qQ��U8�7�j	�a*!OW cj��<����|�aƗyi5�B���SU*/vBԏca������� 2lԄs��P������\��"}��H�--�m��J�;g%�d&��z���RV<[8NB�4f�q3VE���fd>"�X�YoLL���]��,���g��ơ��y?O��<�v�8���⨾��=����BO{�z����b9+V�fi�>7���cô6�-�H9)��(��ˮu��	6BOO,������7��`f�?ִ2�\�R8�`�a%�S����z��A��>'�M��.�G@?\F�d����)=�r�Ț�GJZ���M�|��cJ�}����ɐ#ױ��w�\�7���Y�sؤ(A p�ж�x�ח������S�eu�+}��p��LǊ�u�=�%�J\1�"���e�"wp����@<���נMbݳ���+�Ş$"��u����59U��"K�hm.�u|���?�yp����Oѿ�ĝs�#�M��䶅"��5kkS>q>�A��z�=v�Q7TǦэC�!��PC������i����:�60S��Hg���&7
QVd��u�M?����\#*]�������e��G�ܨ�y�qF�V8�W"�J2�����m<ϙ�A������P�xlL���nN��ߝ���KYQB��`0�ϕ�j�Rh�3̝Dh��O�GSc�T�im?�8p������S>���"qu�W��KAW������4X����611Ah]?}C������#���q:�$��>H�'�)�l���'�q��o�]b�n��W)V�S�9� ��-�CFo�z<�׿&X�����ǔNb9FFF��v����`Ry��C++YhS�4�xpejSP��P���C�g�����PgD1��i�_�P6��e���8n'��9����A�8���Pצ/�{k�y�^���o_<�]�.�0Ƹ9�����
�S��cɺ<W��C/}��s�ڤ/�`i���hjiM/^b���~������%�.Q6&� $�XrO�/Kz��Ǚ�ȧ�S�pf�{�-q�P!��j���Ȳ"�Z��u�j9�2�q��Gtx��F��ň�Y��k^Vx0���n$Ϲ���0ie��J�����o����7�Dn��r�D~� ��Z�~�!E�"u3j�P؂�$���,��}rl�ϝ���sQRW��I� 3�x��lh
	qwCJp�V�#1@���a�@5���M6����kfƫ�֍��P�k�LQ( ᥽�!'�V2`�T#�Bp1�o�i̥����gBw6e���(=C�;��B{���Y��!!	�|
� M���M���Ǿ��,�8D0ӈ�&���52��(Ħ��O��]MM�V����A��V ��^svI��T>yv)��W�[�Ī��ƣ�9)����]ϔ���KƏ�� O)�>+{/f�mDh�$�YiSh{���>̹�̐$Tt�]mh�0��]��z�֯C�X%bYx?���o[��XRh'Ij�u+��x�aִhv���V���:P
BY��܂"��ɗָGOw��J��w^fx�G��Ϋ���g��vL���d��jYV�Rr����.p⸩逾��x]+���+N���l�s��r�pffF(o����Dي���X��;K��d� ``����K z�j6���U�F�(Hu=����<�"�����DZ�M�Y��<�ҵh���_)=1g���5Xq�L����b��0'�pF��������=h�u���%�ܤ !j��B�sleEJ�a}[���{�Ն7.CG"�; ���i�O�ho`���-�
E~"�	�[�����Z�|80%SSS�Dh����0�r�C{�H�����Z�x�_��'�Gސ����fU��ǀ}J��A��
.?�<b�1���ڇavӿq8��ЦXyZS�*���<oT]]��|2����/9�l���'?55Z��H�7������:f��F�����1�+1Lo��}92���������/�&n�IuF��p�o[���sb[��wޒ
no3qފ��K.�=�_��L��@ܥ�"����Rwr*� F�M���N���͕�C	Tht��9εtv��`ro=���ؘ��x����67g��3%¿{M�F����Ni���#6i��4��]~�˅ʀ��C�Μ� 5�D���Z����]������Y��u4ڎ�<@�ͤ��X��O��m��&& F�6T�̏�,�_���
'K���l FJ�J��m��[����!nD�������`��4(1h�	����S�pm���U�^�"& 1kkg1i�eKK���ץ���%����G�o�_��KDz�t+�T��*T%���Fd��3f$�N���=�G@@�n���=?���4 �&%9�\b��ƚג�����2õ����E�Z�0U�yV���#�
"N)7/��0i��2iiup����g�###�{�ȐǦC���bD@����(m`��bt��Ban�!
ms��bA_�豢(W�T���Utz�x���� ?W���x�~=�W��Y�F�����DT㼏�:��^��8>c<ܿ�a&L 귅r�LH�m(D9�n��F;6?V+�"J�,�ԏ�Ӹ
�fMS���hPRʧ��v"��Ԯ�5���X(��;
���\g/"���!@=l�Tm��,8@�4�~qd�����o�E �)�ou$�4��>-�{r��=���7���K�D$�5L`Rq a��Л��+�[��.X�5+''�kkv�6*�w�	� �x�_�<��}���gƒ ��c���'P�.���������}�ǉ�l'd�	yKƱ7���!;��{dfd��!;�^!N�N:���N�w��/}�����8�D�����㺯��19u����t�OO١���C_�,��ÿ��_�Q7������]�E�&m�F�[��Ũ r�/�ˋ�Z|,9�>gĿ�-�e�4�W�,x>ӟ7��lh|dV��A�m�la�d��7�'�D˃'�Z�dR���><�
$ �8jNDR���gk!�{ 
s��� ��
� �ݖ��6*�&?*��;3�n��.���"���V���B��7�t���T;ǡ�<ΠG���>��^�U��k-Df���w}/HD�'G��u�+���[_::.�t*��XYY�����[������G��,>#G��I|ެ�`vv�)Y�D����,jƴ� <���S���[�B��A*�Ss���;Q�{|q�%������G�\Q=������_�>�Hߩs���V�,��'x��f�3�u��Y��N-��،�y�VV�"�痟��Ӵy(;SUj&ydV��o�z���z��2&���2S� B�W+}��Sj�Nɫ����[}������i :��V�b�9#|�hK�ɢ8�ͭo�g�ҫ҂種�6�?�F�ڱ�]����"�W��l聙�L8�TU p��J])�64�����}5�>ԉR2�WK����߿/�8����L��yt��1�#(II��b97�\; �|���R��ɣ��{8�~�-��c��c	��3j��?�n���zn��4�'�=��<1���Jw:�>���~/��u���F:�%.p�M��X���6y�\7�Y�"��ņɨ�O����Uj���@�%i�]��Ij����LU��z�U������l��i�:�r��Kp�J�L�L���#e��/e������̥����E؏m) ���m2����'�8Z*u�Ļ���s��;i�P;�X���q��^_T��X��:L$iկ]Rvf���1$z�O�v��\~-�:9
���7��(ɱ��T0����w�8T�6��uͣ��˽Ġ&�ET9�����p��wehhg�u�[�wS��?�i�W��&�1�4K^��T��.s����HA�� ����v^:��u���v_Q#q^�`�R5���ܺeZg�]����A�NB��[���-��]��F�Q\�t�?-�lUW����M.��g2���_r�q�-e�ܭ`j/�k@�}�[EE��B?���N'~ GߺN����aݩ��]���ގ��n�rt]��SR�n���Y�?n���Ya�-a<pl�j�<���~� -�=�z�)p�,�<����ܹ�x/_�
�ͰT��~�2ުNZ9,��:]������M��;�t��A�\��Rǋc��3E��f�J)�P�A�?4��+�^j=�rA0k����"��Hw����r��
 �����סR�b��}�ʵ�U�Zet!��6D#b����4�XaY7�� h�[~R5 Ғ�+��gۤC;�_7J�����.�"��Fn��|�j�e��k\?�w� ���݊QW�|f ?[<�#�r��fQ���sM{i�$*К��+��q��)[A(�l�h�e�mp��Ղ�����
��_T	$�N��kԶצ������~�$����w�/����@�R�<�F���o$7ɡ^���#�ݹ��gN��g�+��x��]�h	H�Mh�޽�Bp�ɠm"Z�xԿ�BC ,���)�ٜ��a�*Nq��-��ޭ��>�>�@�D͢��$®���i�8� �2�klk�o���¤�+�.A��g�!��N�{�<M���(4Ӂ�?8Q����5�:0�*�S]�
�ϥۅ�vq{�����9�?-d��S}��r]8��I5 w6>�3q�k���sS��\��V��5�4utD���
9J�Z{x�-��n��k'"L��w�<�&\�U�bc R�M��;>��V�u޶O��t$���81�������*J4�4S��I���z���T��բc"��xi�k�W*���ꛘ�I�G�hX��'�2�=%����Q+uZEϭK�Y� �(~�jZv'����$�~�4Z	H"�jc�g��Tq/����1Q��O����Fv�P��o�X�x$7�,S2���Nς'g��w3�gO��?��wiR�����̧�m�=�e}���ݭ.>�K�}J]P�1e���j��n+R���f@}s�Ñ����b�h�������B^�d�<[鄋Y�x�=++%h���"z#�i����S�kO}�S�+��-2av��ٌ����U��LC���ƀ�|�_~��r#^ͮ~z�Ni/�0G!�>(J'���1��8W&
G5���)��ʱSCb��u��U^[K7�).�Jj��- _{��j���rpx!&e0��^��t�˝����C�����W���^ٖ�Y�2��C��YB�)H���h�n�i�8�����)��� ��{���:I�mq),Q.5X��ؘė893�,-wx�tB�� ��K��-e4dLu"?~XX��s��k~����trA#f��+���@�gty��}��F�ۻ)��Pé)���kJ�{5�zz�WV�	��ou���; ���H0����s��k2;�o�o\�9�QR�v�/1ʱ���d�U�	D	���<�ڵt����S:6
�R'���3���C8����[�uG� K���A,�60����(S+����,(��W�їՂ��N�7L��&�<@�5����g����ʃ�)�d��W���v������~��B~���jI���T@:m�G	<h���9*A�O?�oKY\�� ��b�Φ��� =������)�Ù6I�����wD�@���/H�J�^��as�Ȼ�au*A�6�Hŏ;r�w��e���-�+��:Fg������ϴ�����:�����n���Sf/pwK���du7��8�~E�,�%��Q�WW��Y�l���r�W��6ͽ�,�J%�DA�Q=�L�؉ّ�=�3�7Fr�'��a)�p�tZ�EQ$��굎 �����>햀�*��u���"0K�|05�<en�fG�*E�5q���D��^�;��/_��P�>+���m��u�aa���*`�}�ݿ��ktZ�Ŀ9��Gn�������<�7�(�>6��N�	����㱫o���î���^�*̍Ԁ'��9�窕��Kݜ!G��_�;�7��-"B����<:!+Z�F������z��s}��u�G�b��B���2Q	�h|��� ��.aP+�+�C>��V�k�+>_5�t��G!�f_������=$v��j_���-Kr,�R�XS��=,�jo�� �A��+Nt����m�%�K����Z���#�e�����W��}}��u�<{������"Ɩ�����v4� �9	�CCT���:!�߼����x��|6��"z��M����r����\���o;�`Z[���U���u-w�5u�СZ������Q�zu\L����ddG���u�@��|���R���
�j�D�5��g�91{k�/�al�b��U��=�\���[�ɿ`�=dV��cX�K:lO���Z�ë�\ę��yJF-F���c�J��KgQ�r�޽���|���"@���ڦ�U.��������>˗�|󩿜�\��Ȫ�$�(NN֔TK�I�������gF��94�S�,���*tp��aH� Óa��f%S����D���� � �z����T�>R�yc�H%P��2�x��ԥ<�GKKW�L�o΅UO����=|8zmٯ}���~���>����"5�>iT$?�=;�Ɨhk`�s3M#��荋�\_�߄g���w!���8�yQW�1@x
f�K%кs�H�M�,�L��0B�@���ƾz4���]V"[-������ZN��?��W��ϱ7��/v��Y�5]uB0�G�%uk��}����J#~�g�zb�P-�h�gVuf�Wu�˝����W��]-K�z���קD��Qi�U�*^��2MQwq�{�Y8��7	 Ua��)�Y���q�:ec��4y�xC����2�.�Wsg�o��p�w��<}ޢ����}_��~�]M/���ߗ�9 �;}����V���0B�Xڶ���Ȫ��%�Fuq�.#�ި:$�h�ͭ%��rm�v@���2h�BO.�Ǹ[cZ�J���c�+J��,���R4��z�x���Z�U���ܘ��Zgs�s��y���@,�����^�`�kT�7��*X#]�BK��5?��!��y�^�<��;��66�=�"9c����6�S�/�,xڣWˁ_Q@Y[XA��E�H�q�6��O�/�K���%&�k'
�� T�<}���}ꎺ��ܳԄ쩤�ī>��ծ���Sbb$/D�S\,W��s +-��C���tx�{q���0����B]]}Fp�ݥ�\�����A�����6%ԏ���5?�fs���ޣ��r��N�S�����slJN��+)+�c���S��7E�1ˡ�ë����pͳ�r糞�W����Z92{)��*��|�3k�4����NnI��*-Ӈ6A|�2�x���C�w�9t4 x��^�ZK�L�ۊ�n���BOu��x���cƝ>���K�j�&[$��9�g�$6@6r��_��R,R�/�)ȟu����I�-���r�!b�\����v9$4��u8��YK��x:�w����?�rc�������跡㝳r��=�d��LӞO.=�Tz������f�C�E7�����bDa�,��I2!E�yy�Zֳ�$���]����ZZ6�*D�Ti�)DpZn�M�Ն4���>[��g�35%%z�bE���_�D��X �/�.?����Oul�wG����V�b˴�Qg-^R2 a{���0�7x>����P�%8�]�.�}�TI�H�F��HFfze7H��JG����QL���7*��)x�6w���S)��h�Cn��4��u��/:w��ۖ~����,qz?|6�	"�/���:�?�"�9X�uָjo�j mjn����H=<T/�{�"89|��X���\�`N?&'�66o�^�����{rv���MC�etq�:4���8j*j������kJfU�t��d�+vv$����Q0�>7���)j�T���z��r8�'�=NX~@�ⳋ��C&�:ʥD�:՘Ca��e�ߞ����c
}33�@+{���S��찺��tߔ�u��O1]��I��0{/��Ƽ���ΰ���e�_c����'R�8�P��j���洬�&	�Q�`"H�ݯl`��~�A�t�����|,�N�9��r����
������_c.Rlu�/��JӪQQ�}K���{�'���$�����
_P�h��a�ro��}�>���N�CF|�B�� C��{���_�����{�DgM�J��jo�Y�i)|�R�������gi�"� �S�� ����~�פS.R.�8�nϗ�;}�pR�ډ]� �6��2��ӷ�}�"ovy[��e˃�lT0�I�UvAǎ6{3nx���meQ@���z|u�
$��C\���59#�\��V���v4��o���t~�XX*O�fu?x&֦�T �u����q��{U����5�	GZ1
v��Z������{?�[O�Z�O�Ԋ��WY�xO?�?K|��+�����쩼%��Ҥ:���L��Pvvvܛ�_�$����|�stp�����X;�4���&��SbB�bAsݕc�:H��%J��O�V /��S£�|Άhh��ܩ��Q�`��}A�&1�;�S�� ��n�{q�)֫����W���Gn��Ԯ�,�*
���<:!���&5���Ȣ"w�kL*�n?��l�'kN��b���	P+r��}���+G���T8iX|u���C����0^�W�mQ�ńK����Wj�K��_�S0(8{��;A������z�e?S�!���	�H�mmꗗH���xa��k�
$����a�O�S�n�G�ЖC�42�����
����vw;�Fo� SI{��Y*hȈ���4L$��s��6�����^?�ɯG�CC�nn�d���8F��� df�»��6��TӢ	h��3����WW|�V�M�2�h�
�0G�g�}v��7@�H�f8�ƒXu����5&�����~��0��pM������:�P�o8j�$_R�Z�ď�ٽ[߷C�>4����uCq�Ȣ�f��4?������P�ӷ&��4��� FKWs��~M� ��Q�$��ǔ�=�����w�3�Rq����(V}��������e�ݖ�DW7�����+���%��^�Q^p�u����� -b���`(҈�K0� S�q�b.��V<4^�m�5s����ݒ/B���R�܀7�}W|����f|��r'�8%��[�Q�xj��_���䚟����U7u+�����1V0���%zJ[z���Ŭ�������%���72V�R�1/�恊��h��*�X���{����7���ei-!�4x@`�0&��qSpg<�X�m���l_^^��:��)�m��Z�f�2� ��!�פJuA-��įr14���q� )A��'"�駏�X#j�f�[Yyx�\���������<�^{~�ͣ��^W�Y�Dy�O??;�6����H���WV���]��i.HO�������C�nğ�[ѿ��ܪn��#,ybb���x��� D��ښ�A�=]{F�D��A澎	��}2��~�S�4�d:<!��G߄×έwoO���QwZqTU)c?�L��J�kF�/����Vl���u��[�isb^�W[ٙ��tQ���xd����wԻ�c�~�-�SQ�W�4�^�yP�~|i�,�d����Ç��$�z�a��}?W�s��@�����������COKC�.8�(�����r;I2��G5����+i�_���СB��M�3��1�jC�-��T|�����<c��ub���hۆ��Yw���U8;\W���}BPv����>����O/cX�gi]�e%�r�
��TІ���_19��şs��EE����9:�����ܭӕ�Jc�0�ㄑsӐ�'Y����
"`^?���Z3�P��q�uڬ||���d���}�������B��~|�d�R�Y����K����)4ӹ0[�u��cʝ��rB�~�ܿM�&����ӈ>}{]��jGH�X��~<g���$N����p̱L�"^h\(r��.�>>�V��}����޿��i��  �Q"�������~!h'�E颔���? L'&|18�����K.ͽ*�H���m�3Ĕ��p+<?����Z|����͢J��8�4(^&��XI�'���n	�ɉ֫��e�v�HI��yJ]�j�9ƞ�^ljZLӀU��ivy�W��|���nbbr�5'��֯�L��a"��Vj����
|k �ۏaC�J�ll�����J��K��;�d*���Sr�
�|df]:�d:�t[Ƅ(^M��S�Q~Ƌ�%��x�3�K�_�d��Ƿ�?9eeK%���k�[ZOR$���ʮ`�z����ܣ�q�}��F mўA�*rZC��0$ �}S�t��=.��ĠN��5�O
X��W��ńI�=���7��i�ԃ���d<���3い ���w(ܸw�{�k������'Ζ��J%O�_?��e���P���N��'�Ǧ ���;���s��)�5Ga���*%��_��&�n�o]����@����Ss%~O�Þ`����0�5�`����}������*y�Z@Aǝ�z$\��h�hƞ�����H�\cˆ�ʵY�����=�f.�10�2==�h������h#�;������s�� W2ȉ ��gŌ�U��FʱӄP��3�����?N��{b8����h����"��:\���'���K���ޣ�ɡf� ��DS�
�T�L�8�˾������ʉ*��Z�ZUZzzay�8όh��aUX8{�C@h�\�/�KX��d�y��֡,�//��V
U`����k�ȽR�Oy,^W|\MD]gU4?Z ��ш���0?�B������!
�|�O�?�3����s����j[, ��,w�uTK��~T:�.,D:D��>��{3��x[WWW���]�Hp����+yw;M�MX���M�6�!v��������5�Gɴ�Z$0�Yv�j[��/V$2�G������ou+�Lk���
c:�`���wØŦ0���}�߹��R'�s9��y�dnJ,��a��fya�@����O�l`�H��w�:4���o���jL��d;�}tp�>�lf�L���MW;B�!&�=�٧��$&|�@�{�*ll<�Я�4���7Wwq��.p1u�����4vh�h��#x����R0�����?��i�:;_r�>���;>~atp��*Ū�B���/+�,����,��\�Ƅ>.�T�:7���y��E�g��J:������^*j�����V�d�ĳ"��8�4��ğb�w7�������1|�ňpwI*qx0��H4��mӅHfJݴ�h&�[�_��bۆR���7T:!ae�MM��GG��~���SY?��B"��]NE�	Q� kz�g{yn�x�)��uV�:�YYE
�����'_�$�'����o������J�0KQC��S��'�ŭ�'~WcS���K��q��r�Bu���x�:?02��7l[G��'P�`�=��&��ER`0�ջ�H#22���MS�;8;O��z6/�&cK�%r�˙׿����i���̅,���!R�4��� }K;���`�h����
�\� *mr�� �?�������J��!��r1 o�ӷܴ���_G�
8�o�u-|���KsB�D�	�ҹu��_��ς9Ec�d������b��jL�;O.��N?I���y����?=����n �]��r��$�g��g��z��Bv5jz�m��G�$��]�4��+�͋�z	�i�?r���7*������N/� ��T�ٹ��������z=����ٻW�|Y���#�	��O�5�x�c��3H�!�;B�v]�Qa����~�r�tx�K���}�:߸�E�np��3���iR�q�� J0Z�+o{�|.��35�O�SO�������22qn�Q-v@�:2I��i�����s��s����~�����Ch�=%�Wl��Ӿ������}���2=�?�u(�>1��k0�%L�O����;  ��z��F�P���j�����C�8�XHq{�>���3��qtU��Y8��+��+�A'��	��켼.m|WK�,yKJK��>Y�B�ዟ{�\� ��$�Ǎ-������7N	L��[�6K�`�;�Q��f2�6`	ع���v����A����t��a�/Hٱ��D=$ҧ�:�5���wP�8���̫�;�����|llF-Q���ǝ��C_��������6�.$OF����OQ,�u\����'�j�ܱKKW�mm�r��smv��2?H�w�t]�ʛ/�F�6�DC����?�z�iIu���"��Y(����/Q[��5��n���?ݔ/�H,qsbMg���u��Qৼ��-�(�ߥ���%7Imxq�{u]W��"T�������6�4uݧR!��Ζ�-saD:���/_��N����y�Ŀ��=4�S��|{��[X�Rb�/���C�����A�|'S��#���Pg�W�-mZ�U��AKO$�5s2�V7�-d�Ȁ��2��j�����32<�I������E^���!��HN<�;ې���)ڤ�d�e*3)ָz����1�dQ���00���:��Pewh�B�Y@�r1QP�2�e746&:!KKUt�3�+a(Nt�ǘ�V��a�,
D4�(���r01��5@�]Q���G�`zh�������%vY|0�{�-��r�EE��p�%���0��B?{Aף;O����W3ݪ�j�'tr?��z�5���F<�"t�ϫq"X7�4�
��o���K�.�z{I$�@��k���i�qT�k�d�������.�,�̼2��#]�?��3Y�ך,��I�}�[�3�����ۆ��βm�R2���MH;lu��Ӗ
y,_���8��U@��̀��@�Zu�������H��/�n}n�3Z�{��-G��Ӳ�xJ���Nx�Ë�����R��Pq4�~.'YnQ���넣�Qʽ}-ҟ�i�v�W�{H�#�����S�9e�h�VE�7����!]4��WjUW�]���mc���Ã.w]g�"��|дF�ږ���$"�,M8��S5�/|����s�������,����������_��B��@N���]����RJ�U�m(^�.`���~��߷�/_88 ����=�G�6�:
}�Ԧ_��-��e��I��&$'���5�_��BZ/��H�ۦKG� ��Wp����������� =$ٷ�N'��%���.0]�I�_�NOp�0�S��`X~�2�K/Thhͤ�B)��:����S��3�}1��t��vK���(�R�e�#��_[@m�~Ӯh��\����nE��+��/��Tܻ�?g+F��������N�t:����g��\(��/_h)b\�O�:>�ڡ����V`_�C�3��k?��o��ND���q�;<�ֱ�F��ڞ+�irF��z��ˬ��E�cL~)�y��	\���d@Viy`��p��=<E�b���j�}-<��e�o�/X� ���Z�E�fK�y7�p�j2��@H��
��>�rQ��>R�#��� �J�����`]�d]�U����m�*�+22n0��:�Ak�E��,�t~c����;kp0`�)�ŗ�" �hk�Jd8��2�zZ:e䦡V���Ȱ���0��+߲�<��S��w��P	��� Hem���/?������cY�Ŋ��o
Z����$t�,�,��YF\�m�I�A#�	�F�N��@?��*~�9ְ�Q�ӊ����K�:oi��]e�9��إ�zYFzK?~ժ��P��T����OO��+]ⷋ��F׵! n�rI�����M��M� �B�xjE��?������yp�uj7�blo�~��A�K2��	�̶�fW���cCS����L5�:����D��P�(E��c�:�y Ю�+ a�%>�M7�����>p��oi�ll쮭�#��$�		>���>��uK�Q�k�[�����/Q��7;e��l�V��D(WU�-
3��n��p�ĕ8�/ٿ��{���/6u�yU(�a�G��կ{X���?+��2�=�yT�;%�s�g�������Q�l�h���y��4�2&��u G���O{y����]y|�ͣ[�z`lx�8bi��SvV��ux8uY��#}曚������ͳ(;����ƿc����}yy�d�l�dS*+���n�����@�9��}�:Q�bu4���:���YC����`�(&�cWC��~u�A�����9��_<v��g�*קIV[�n%�򮑢_H�f��ߍ�u�R'2`z�k�M�}�LBU�
p�R���|� i^�(}��|�`θ�8m2�+2@nTF��2V�9%>��f�[u�a���Jm��?~0�'��@�鍩�E�{�_����{�H���-�x�d�ɩ�^��k�r�� �����q2�n�Q���NP�3Q���=���\������u-��
�n�g���O@PS�q\TA"lA����|(]��ӭh2k��Yt�	#G�󁙝�M�7�1y��Փ�w�Ybs��H@X]�8�7��Լ�[,��{6��U<ֻ�ݿ�Iq"�:}�$b��0H�k�;���G������};6�F��n^/���Y���ZY�r�S�wii�&/���ŅYT�)�0�rɓ.ZJ���F� 
(��.�߆�g+����f?�j����jɓ����6�͗�A�[t�
�u4ԿM6��Q�?:z�Ё�"p�0�:�Ѝ?��� O�"2�("Wb�~qd��˖���+D�ȧ;\�/N�8̭��1<�͍�]�-�x7c�z�<���%�L��
�:��$k$_���.Lx�$��| -��u�s�
KH��V������m��WdW����y��\Q��M&a���8J�M�l�E�;P���j['��;���O� R|}Gw�j���1���<ׂ�X�H�+�ǬhU`B�hT7��c7��χ���PH����:.����W���Ī�����869ۉTM��j�[Ȳu��<�V9��5��`�S�.[�n�-�������(@�F:���&=��¶K��tqpɢ3
��)��c����Vu�'�889e���r�>��
��� ���2"A`aQ�8Q�eD� f�k�c`|������e}�r����%�I�0:��A��&0�|�2J���zrk�^<{c���@�P�����
��I�i���[�Ӝ0E�]�x��7�*ol���H���:E4e��0�IG���+A9 ���o���b�����`ۀ;piN��P:/׀�
m���O�?�p.��R#���B��ľ��*�xW)�T E�4Ҫ.�	�]�Ks3%�B�x�M�װ�S��!5a�P�J���Q�p'T2 忬����;M>�'I�_����FSS���j��Ys�/v9 *��S<�?��	K�k�����;�Z��|�q���J:H\�#:��U��d@b� F��ʮ��T�U܂5*?~	͇�sB��;�P�tNq�]�N��n����Pͳ_���D"��`Fj�d� �ƅ�^NA��T <ew<[-^�T���ڹTB^��P�.b
? ?��q_���˃(1�j��S��r�:P�AA����`99��pn�T�[����_>��i7�_��7�ɮ�����[�����x?�`q���'����g͵�p��A|����T� Y�,]^���_����v��?n#�9hP�7y~�����i�Akc���|>
>�1��N��Z�Գ?�0�~:�\�?~���:�rr'�l���!`�s��voTq4��.~�;�npv�e���~���W`ң�C7�\&�2��l�k�_m����|;�R�� ��e���9E�S�P@����xx���Pß?#,�_��\�rܑ. ��A���^.�e8ޟ�yu�v�	���g�Q�lEm�4��o��BL�JN"����(��T7qW;��L��*.֔�/���+m)�(���ON�3����y�-�,�l�~D��* �UW��ҭx�2��ޛ�=�q7(~mT���ƏaC�Նjh����#����=�s���י.`��y�#Α�$�������}�!�v)B<��>Z 166��C&�3�Ō�ny��s���T�`xQ!�%��sO��Gǵ՞ѳ�A��[�]�@���9ܟ�����D�+q�a*�A�yM���%�l�/o,P;�rfJ���
�����B�Թ�u��a�� #X�]���6�-�g��QGy�|���c��J�Ұ�!��Yں�7gm��S�C{{~㨇#*QQ�������c������NDO�'����g�׬��C',�?�n@������^[��$�[��]�����"wi�rN����"j=��~�����nF��^�#w��e�S�Z�9]����}��Ҧܺx)�_6B���=Ju� ࢋ��q�]�B�r)w*�Y\�������5q��-.m���-w�cS�%����Z�x,į��^���LG����(
�s� �!�!d��j�h��&"#WYyӆ���B�v5��36w+�Ɇ��l�˔��K�|Q��6J@�(���/G#�;ǝ��)�e@2:�A����	rb0h�u|��=�WD�Fi����	��}hΤz����:�/q#��bJ�:df��U�t��	��Ŗi�٧LA]~!�2�W�f��}#��w*a���.��>E���L��(`f���.�	@�����V�Ւ��a����s@n����#�`��)-t��v�+yfff�9,5�F#�u�������߹߿.��vgee%�'�DC���´,�I2�8<ԓ�����vφ�5 .�G�Ã�r�s9Kܿv(�B�k��_�
�\>�6hAL���Vi�uǱfhQ�}V�i���P����Z|<��C�� u�H�F���MK��zz�b����]�ȒH�G����`��
],`w�p�r�H�x�ٷH
�{@���ׇ�4��}�|�<��d���\�P*_\��[渀]�w�ýϵ��{(,34u{����r�Ç�(u�ȥ�+X.hOf�cF�n
s��8#c�{������g�SR<��&���X<�`��nf���QۆK�Eѷ�uZA�҅A*�,Aio_	�RA*B�/����1�F���#e�s�%�+��m�
V	�Ԕ�uM����Y"A��x��0�31��5&�K�Ԫ�T��]_T�7�%(`_���5������$��JRZ:���M�S���������ͯLOߚ$U'�� 
�9	(����l���d�;	��~���vV�uJ���`B<;{&fu5����:s��\�O����C���l���E�/?^�+�Ʃ$v�VCok���Hrt�V�6�w \�q,t�Pv'-Y�_�}6�?��"��Kwɨ��8��g�	���аn����V}@�~�S�H� qy��p�kg��˃��`[�J��wyu�M��7�|�\^�r�u��P0��R��H��+�ϝ̥
wc#�k!{s���d��!���_�ږ>� ꥒ�jS�񃆴z�S��4�*���}�h�d�j�3g�J�$�����5?���z��K���.S�I�74A��j���_:��t�*U��g����n�����s0�G�l�����I��LD;��Y�x�M�����_���'�&�/Dr�.L�BL���i���ݒ�Ḧ8���IEI�Y�����[�7+$?��]���
'������m]s�|h�Ii�
@�, xcbx�ŀ}𠠸X�3M�����r������ /S�s��Z:�i(��ԡ�%�z��vz�h�@�n��s��	�rR�8A��@��ܢ�K��tt��#$�d�k*��˯��zBo�� K��'��������ᓱ�͏�>�Ք�?�pzfU�p�j��gF+�{N��5�s���+M�>�"�!|*��-�}���t���Q~�! �}��Ŷ��s��-�������x�����17�K\���ǌ���{c�9���1Tض����
 ����\�ڶ�v ���G��T�a�yaϪ��uɉ֤9ޅ�E7�.h�ŋ��Y�k�^��d�iEmUG-_�a�ܿ 8xi�6	��' r�xH7R@''eB�b� ��!��n�],��_�v	W�ԡE7�����=-�y�'�?DOׯ�x"�B2��V�,T�X�,��ӻƼL/�a�SҐK�y��ʷ�Mj �����	��d�rs�krz�)}��ٙ�Wg5��=^�W�U��
:��)����<M;�l���7���������Ҳ;��A�P��_Kl�?HU���s���`
"*��h�ZD�;�����B���o�y6LN�W0�>��4YZ1�EC�V������μ�T�.�[?���� ���ڠR5 �㮥���E�����^���>�r؍ ��>��ù��*�����v��q��:����RRj�s�1�|p��x����n���saooR;8@��.%`w�W�'�Z�,wҲ9��c���e:D.��m|}g}���Qg#�+!�n"?�q������U#ߍ��0���Sq5����?թ���v�yo�iUU��F�����Ֆ�,�rn��f{3�z\��,�<
�o�b畩'ں��� UlӒ���@~��Q�eo	A]TBr�A'*6UNf>���"m��HT��9xz���ei��~6�sH�Q��..䮮,`�Qm��]G�ބ��g)�e��U��x$Ze��<��"��ٖտ��:^sњ�Jg�_��8��:z�����>��{�z�����Z�-�c�4���+��y����	���,�LH�����ɿ��e���/?�I[��@�HgIҐq�*b%ž� ����nD�T`/���h��"W5�r�% %�NI�8�/��|l������H�x *�2[Iֆ���{3�~^�>����ȸ�#�SG�s�ŷ ,����ڒ�V�_����Z�X�p�7`'gB��TC�����l�������Vuvqc빀�[d3?�w뛚F�� Q6@������@�oj�st�$U�ht�����a�����7�@ܼ�_�8盤�Wיbm:���]i�R���R'��&"�0�gb���E�\BC~Q����H��@����g�����4�����;�����h^z�`tٝ.��+UU��c%Vu���=�>�V6�$� yn�t¶dw����/f��=%Q �����۹�o�zl՘���K(��{!�
���d����c���B���ݵ�;�nA=m,��T{%|3���/��P�j�~�Lv��݌G�}��r�1�x��P\�.��B�0T�L�'XF<�����N��p�j�p�=jѴN���'A�s��iu���n�^�I��r�[�����8�b��Z(0H��ބ��.x>��9j��Gk���E1�Z��بH��#�u��m�����A����.�bUd#1K]��b:���N�ͩ4�T?��=������FH�+ ��ۛ��{�|�Db��g�H!%<oG߭p����ݐ�������v9)M۬����}�^��eil��wVV��9���v�!hr*��,��'�3�8�0Q~��-�x��o����{�yM,�pm��K�J��N�7i-,Ĕ��=s瞧"���˖i���U ���f�S�,l�1��r�P�OF#�[(�GG��U����jsѐ��_<̿NK;շ�mc�p��1ć�bx��`��UFǂ_�'��[����0�����
�-=��_���tSZ	ݓ�ut��|yQ�����1Zn�ST?x,t�/�V?$_�``�8��Y���&�����Qq����
fhq���J��c��O��:~V��G���hR�tX��ة<ՑXċ*� 2B��!莅���! �/L��-,D�����*6��x�~!ۆ��&V�8���m0�F�D�'T�8�J#}>��f�@gX"�*-w���hhC��v��?<T7��Rb����w���J�֭� �bX���A�����b@��b*Wāg� �`)���PV�L������bz8c��۶A�����k�(OJ*5�8㩣7��/=X4�����V\����M��A��U��a� ���S�Ҫ�1��ٜ���_���s>J`x��� �Ȉ��Óv�C7�t����!X���.>/F�����%<����	��������I �� ʰp땄2��"'��ϟa�̔�m���9��B22qYYƏ���\���ڡ�K�eV�jA�<<����#���2;?~0y�=���o������ˍ�(`��a�,��$����D3��������=7���0�FH��R�g��,R�X��2��F�N\[�6�ilϥ���6p�Q(� ���\bR��g�G���8����N�J�_��{�>sf>�x��>�IT[9tt�>Y��Lm��S~�2W�>E˴�x<�$�Ѐ�H�_>�@���a�Cm��M���|6bnP1��_�F�qc��i�4������3���{�P�}	ٷ�$�dߍ5��dI�}��}��3B!��&��i��������������?Ǚ�o	s?��~^�{�{��F9�a�H���u2�n�zuȝ�����U��!r����{���O��/E�mks�7R18��+9fO��wփ�3G�}8�'v�Ν���V��r�ߤ��0-�2��*l�C��DO�������v������y��,��Q !{@�~.��g�yb:#l��~N�����м<��*sL���Je@g�7(#B�d�z�2���m)A����R��$.�P"45?�<i_IA�R� �
��~$"�\艡Ӟ�g���g�8�6b�F+��svv>n`�R(�����x~��fF~`�����6���J��M��55*d=��/�F�D^�����s���J�X���߶>�x������.�P��6.��2���Vю�Aq�#�F��t�����$~�e���,z^a���� �;4���`�̀��E��y3Q���+> ���4��NN&r�������P��.CZvq�ؠ���m��t�f�	W��FQtϸo��.ҭ6��ܙ�(l�.��0Ct	����4_G~�OYOD�)��AL�?(�&���C;}������㬷��ʚ}��{Rg���*��|����%XN莬��s����!~� ��Z��';l��7�5�9���5l��Jx��C�5F�):��J����?�\�����nDP�Y�3o7P$�e&63�HquG��
=���*U�(�.cx����k΢�a��_�$+G/��zR�d鬙�[�5``�M�\�ɕJ�W�����2Sd]�6�r���8b	�ե�8	8I�zJ&�zQX��Ǫ��t.@�Ӯ�\�y�W)V�4��������_V%�kl�R+z�w_Z[;�YM�[)j	N����O�l��q��������u��(t8\��ICE�址�?G��x	� ��l�C���Tc@̭e��}К�Tf$���q2'	ȣ�Ww���,"��2o�^��U3@AxiՇI���bH,�p�ͦ_�Y���N�S��G�����k/*[�P�va�a٨?~Yt�r���QHP��+^�	'�a񣄸e.q� ?����8Ջ|�*1��P����S�κ=�:w� ���h׮1�9?���CF1������0��+Ɛn�*+���M�(0���<���/��X�Kр�U���<��f֥?m��-��)&��� �hI�*or0��2C^4����M���q҅*W�|�!��ƫc��J�'*z)"L��$�dAZ��r�z�x�W�h�kKB{�-����,B8���ip���G� �dέ�v�@�cn^�q����ߍM��T�Ѥ��|��F�H[*�L��ϗ�Ӗ��wrm̅��nI1j��>��{�Ui����iu�<e	<
(����qޛ`�t�3�0"`V�֨�[*ՆH���ۼ����v���?oA���X��K���hdT��s:R�Y�m5��^���Q;�HP�&�e����&����(O�,:���I�����|l����Aލ^	�pF��+�-��|�7S\�hre��'����&>��=�b�a�o|���fl�)��#8�̭ˇ{��KK�7���x,��������c 9������#w�)����\/��0�M��o왛����;����L���S}ڝ bQk�8
�*�V��Sy���&�ه:�%���cs��N�"8�����@�WZ�aϔ=��q������rne��r_���mf��,���JW��٨d�
�����+���r��_�=�]W���p�_��H���E�m�O���͸w����i��͍���5;�Qndj�(�ļ�g���9?�u���d�y��W�B�������[&������H�P)KS�u|,(�E��n��ŝ��Tq#�(���T�Y�g��˖�J�~�Pv�+v���&�28Iڀ�����������1>Q2���I��lF�vg�e�g��/��C���& (]?A�bۯY��(����9<ޠ�V�B�}
�PA�H^c��M?�/�.�}z}ʨa����U�?G!�O��r|[�������J�����x��B0L�>ց��O7��~}Ɗ�=M������*����k�V��I¬eB��L
O�d�g��j����f�&fW�L�0��V��|Iq���]�C2�3<��щ�F���I�?z�_f��=U�����F��Gls?�{ʍ��|�:1�[_��|:��?�&K&���f��$�sa����ki���AU��l�}@̬ll��	!k>�..=���"o{z��x���eX}9�n4����ا��NK���b<^<?�y�!\�Il�|��5Qze�[Nɰ������F�V~��GG+���xI��ˋw��:�_i�7\U��M�d���2����3R��6��:����n��b�Q\���2����<3ޘ=�R=��,n�UO��9�~����% ���

]�G�G4�7$���1+|�ӝO����ϡ�n��?X^]MG�r�s�Tg��^eX��鍻���Dn2�_Xș���� EEDF0O9��vv.;4�>IF�B��wxb�L�� ��  �'����F)hg��,�.mX�z!��I�4N���_*ֻV���L�ĸ4��%�Y�����~�O��{-%>�d7qB �n�n����̔G����yw�rM��Q�H��*��ȝ�*�'Ԓ��{�N������';���߼����ki-|K7SX�9,-���5�qz�f���j��L����ןk|����,��#^��6UcA�U�{p��������8_�bI��x�q����Ĭ'{!E�:BO���h������X�;ifh�T�^P���r-@�`R�0@�����P� 
E��A�:*`W�f݈�����������q14L�~��K�v�mr�����@5k�A���k�L���U�?{��O�\��ӧO�i�:�7�^W�E``*��о��q0��7���5��G^�R4��]~���<M��=�v*���|�.�n$�p[����ёn©5�8�֭[��ƝD����<��<��YYY�r���c�P�uq9Ǟ�_�d R1N�H������CA]�цx����8��gN��/�S0!�OL��N�
֑��#O�����֠Ő�S����ư�z���Iɨk���k><y��/�$u+2g=Z��M\���߶�c���w��)�w%S�u*r�iK�/��]S�u��4���pټ�Qh<[k�l}�����8®;i��2M��~�4rdD��,	\�hN�ʰ
:����C pN`�hI��vt�C�	^W&��hGt]L�Ҽ�~��gda��0��x0����ٸ'Z�S}���^f����z����D�Ѥ���K)>�.(����㮆����
���T����م��c�i@��	d��[�7��~5l������)��-
�01k��'<�Ȉ�i�W�K�Ҋ���O
-Ԕ������XԒ'�n���O G���Rl�g $4,�O�@�_����_�*�#` Ύ�4�#W5���[[%�R���U��
*T�fv�%�_��/w����{��� >Ç1v#��Im7h�[�J���%ǯ����PV��]ҫ��[[[s��cO罂.���5�?1311�m� ��p�� @eKKO�����Z2�(A;�S�ƈ�Z�w��m[�v���NQuړ+�/u`�/�B*�k���8��㓗:��4�'�����-��!/ߤ��(M
����z�㔥�FX�o7�T3��@�_Ph�'s�%�!�om��Dc�@�C��ǫCv���a�{��`p��f-�CI))���M��Xz���p�v�rr�"�K�P7x�����p}/��5�����A|S�",��W�Kn�r5����)�r#��������`f7-q!`'i�LAwx a:k��o��C�i��L��l����z��S�pT_�����0>9��,n�߃V��2��S��3�=�f6by�M�o�ђ��MW��U�B���F����w&7L-,���
й��4{�w����t��YnKQ)q����ܦ��@}�ucB�-4�i�E�z�����CQ�^O�A)��	�ؼ��$5ogIiZ�~���J�*$$�t��U�cwwR����Ζ����ww��p�}����c���12q.�uΣUXT�Ġ]@F$����as�T�F�W�H�)��:	~2�B� �'��i\".�+���ٓ+�n{w#8�o���MO&$�*2�L�W���n>�!�[Vl${B[�<�U�|Z�5BQmH�DYg4���Y5���(�&ի�0}eѼ�m���C�rq�̀NP�%eȁ����In�\𰴱����b�r%zw\)w𽥯/##����իm��m--Q z7��P�FFʠ�������/-1 ����1� �A	��V��3�P}����� q_{�xf|\L�* �@6���ai�y�s@�}�3�W�3�$G�+�=�����9�	v�'>-2��eF�D^�.)?{b�K�R���~Y�U����JMtag'i�zkϲ� � 
I�"��� 	!(��d��N���̔���OL\�7�F/m�m�.}�O�I�FI��3���񀬜����PY��r��-���
iS3t���������������SV)��A�i߿ߖ���I"6�d�D-[9����Q��[�u7i,�������mb AP
ޑ�� A��5��/(p�����U��qe����/{����PFb1���s?á�3��逪?B3�ܚ�q���E�@΀a��� �dSK,ȭ�ͨA�YB�I���N�JI
0�~�.�q���4D����l�.��7��GC�5�构�zɏ.o=�>@����R�	~��s7���_�9�i ��Q�6�Wid�\����нw|R��:ghk�$0��@&=T^Mhj�$1s�f` � %Hv|��WfN�o�:��qc�8P��O*�\*��%<1�zh�-��K/((���摲������O
JJװ��l{���X�����P��M_6���o~V�H����B�9t��N tѹ��R��,^�z��Eo P E���׫�dA �ܞ�j�0��C�S�����q�ěb���2{�A ��L
���>uj��;L�l�n���?ܪ�����N@w%�h{�%l.֔�"���Qc:������TT\��X�U�	���m���<�e�fw%�I������JL�c (��M�@�ʿsA�=����婱�@����(���V�M---�zx����� %�Qkj�6��)����۶��U?��d��ٌ4�yAS7�ɑ◕7g�j��Ah��]����X_w������EՈu*l�%��efC<}�"�����:��w���Ia�DYY�/PlX�����/����*�檝澜\2���|���e._���Ù����@�\�Y*�TV�f��{-GLx��c�/f�_�ǵ�߉A�[[�X[D-�:������	ڧk�[�N.5[����屛�+w��x���[^��Z_ y`@��;6�"�9���P��X�i�����޹�^�Δ[:��ikO?�C�2������3a��U?�*�,�r���܆�Ā�M��ųC,J�T���л����}�����_�R��J�)�G]�N#�'q~��G\�<���ee�j�Q���@فcR*�y?1qh����4;��q���91��S!���Ԙ���j屷dd�US�y�/�d�;4&4�[��� ���=pۮ��d�x,p�X{����OBg'S����+#�������	,VA4��ZV�|��bMq5H6��D)VSKC|��,ѭ�4��u��'{��I��.�%L�֚<ƨCo=��E8�����gD�Jc+'�)�^�6���T�繆B�\(׮��ރW��ȃ�TF�LS��� +�T(�m��q���˓1 ���V1e5Y�x�)���Y�����,	�q�:͑��+)!��%}��<?ur�����Ⱦkn�A,A�7���keee4��������P�4\aec�9�ǣ_uYȎW@���P�ںW�}�����v_�v�$���1o[ZF0�z�Ӭ�GG� -�т�u�ϣ޾>I�X�Aw<���&gc��� ��(����?�(Y�Ir�l�ԟ H	���NQ��bQ�wɑ��٧�|�ɒz�p,7@<Cΐ|�w)�S5�TT�:����/�˃~�z��I9���À����A>WU]��6'&�+�3M>]=������ ,[Z�c���׳��>�
�W�.|�����	��|�DG� �
���nI�;H���Y�
ޱ� �k4����oq�D5������/��lF��7n����y��;�oT{�T�;:"��weUS��ۜ�g����յؤZ�Y�l?�����5D�Ԕ3�z�z44I�Z^�Q.����hdUu3O{���7t�	�Uڳӱ���q�����33����9����Ch�i��[eƜD9Q����V�E߼٢١j��J �m�v!�>�����?}X02S+Y�1���w�)(���=�1�����/.�WQQ���g�$�;h�������ttt 7z?}��A%�	i�c��\�ʾ^b$� $��n�}�10���b����Fbe�}��:�%*] 5@
_��d���oX'�'�~?G�b���֖���G�9����&&`OeN� ������L}�ߏ@�3_Dw��앍�N�´�C�`�>/���s&
'�(��+|�/��~�����>i�J	G�zhJg� @�Fi��ç}^�L�n[���:B�:��4��Όb�I11����z�£�r�vP?���������/z����˗���oyv"��e��H��-�����ݟ��8�U5���W������=E%�l�?xfׯ_oJ,	�FYY[�U30L�' ����ٹT
�Z��k�Yu��9IEwVY>}JVf/���%�ܛ�����Y�����4N66oJ�����nY`hN��'�t�z���<{"Q,�?�R���,�"�,���25͗���E�hej\%��z$���'�G9/5L��J���Z\g���$?/�|"�2�tc��Ia6&L�7B��n��}i����)iz�H!���$��o�K��_��/�p����8�:"�t'J�K-=�?�ɒ	D����{��/Ez��g��-7����9ڟ�f()��蟞fO��qE=N�<��GX;��MM��v���;u��
{�������T���]ts���ѭP��v��\�E�֭���a��l�&�{	ż���
+���&��{D�9�nf�y�k�s�en�,L�E��3�S���s�b��{Xl�,pY��Ҥs��.m��)!A�}�
p�غO\��h�;�M��Õ�� �;��+��Y��L 9��u@t˔P�����ם	�8� &$��>R��s|=|DB���R8���cMMMnVJ����
�����6��n�޽S5�ˉ>6<E��5А�Xd�����������7=�GX�ˎ�U��3�*��²�.�|���
)�;E%$�m<>՗�tuI����G�(�0�b[*�x��,��8ċQ��T�$e��fg�H�p�^�a��a+�74��PIR���2e������g��
Nj�K.	�*֠�t�N����1^�)/ϝ&�h� ���ŻȒ���+��󶈳v�ۊ�r��y��˗z?��Xs4/���Ϸ6\������-�mv����ۤ�laЀ;�\.�п�'^V�TXR2Fg�%A���������,�O�;�
=ۧ�G�w~}TЙ�W�qw,����#B�[8�M��8汱1�ZO.��K�����|����Ǟ��E�@a11���vO�&��Ǳ�����p8��A"SCm���	�H�*�~�S�)�@���ރ��f����D���+N����q���w�`��U�w�N~��f���gY�Wp��>B�B?锉��Gwg��̠�S^��<)��~�hӉ��09H�_�6��uv�N)�����<�<��k2�٨���K�A)dN�k'Y�� u�`oY�����x�_��l��1�H]������Q������|�DP֭��������e�iS�n��574$��<��jo�����e�Y1sXz�W�	S�Mm$5�T4�BЬ��RH7pV;S=6���'{p=��q��(���b�C�u�D�g'��I�Ɨ�i���?����^�K���<�0� �c�u:��& '��T�4��i�����EyʏV�I��<��
��v&y���/mA��w��}� �QH�ڻ�-�'��S�~���\J��}��	�̈�ժ�"�AG �k�K�q����4y��[=}��8��]���(�}m�����]�ٍF�����x����A���_º��$��RЌ��`h�D���� ��O�pI����$^�*��R[x1�7z5=2V��v�O�f��<�8D��������K�dsц'��4��>�u��[�w����쪪{~���J������V�r�!��v*��Q0�P��7�F-�O�%V��L�����~/H6fXի�śW�
&66hrds��ʇ���QP��67'BW�9t��̸�O���V�3��N�4�56�WU��cJ
���o��I���ww�+�	v	
",)�n�ޘ����&��� x��)��?�K����ۺ�ip^������������ʺ'm58�[�]6��k��P.�!`]b���D�z'��b^6��,o Q���A	N�$127�s�Ӣst���F��'=~Z�aX=^�n�/�����[-k�������D�\i�\!��:���&%kS�����&ʲE���R��3�p_��&7�F�������?�:͕�2zvv.�V ��UnII�V�Z�:\~��N���"9)������a�/,���	���{������ҫ�kl4��J������lp#U�$͘��mr�C�лP��A>���6���"�cx��Z�OkclH��{�\�deto��`}kկ-h�C]7���9yvu5=c���=3*`ht�{��� <���QB١1�Hp���'�<7�j�NT�{���M�a��Lh"x7P<<�3���в�X`�"�6�S����U�WQ9#�5�c��8)�aHD�v��3}@�1��
�e�J��ױ�#>��!׳��f-�g�h L��XW�_�s�β��ols����̱�v��q߷o	k;a�/0�hy®k�.G:j\\��o\��>�1$b��uo����3gPU�l��?DyvPv�}o�%S��ۮC�yW�4��Yݛ�ݘ��ȝ��X�����i([|��|�d��e��@,(I�߻�']���/EK�$���� �_0f�Lɔ󵇎8����e��-I�<�m8�"�J����L�ͮEG.z�wWwL�
!�_����ʘ�}����i����_$�HS�
	).����xK7������ʼ��yt8F�7���S&�ir�v���7  ��i0���z��B���W�R��)P��r��'t�̅�x?� ��-�w�V���8�����!V��3r�r�k�@
�'.��0��b���0���DDl��1k>��2e8f�+8Q�Z�w���n� f&��߅�M�(=���(��$"��b���IS֎_T�~Y)`!�UK����O����}�f�Ď���b�2Q��p�	��a��k�ݶ�A�u�OwyL@2���EQ�4��>@?��|�ዏWOJ1��%�ݘ����C8�fi �<���_I,O���Ɉ�?�
���3��|�+�ZΆ�����W�>)����
=^���0<�NT/��k/��9B�΍:��o�C�¨���@���!�Q�Pj]�,����D`0?���2�弲�ȝ\q���q�����@
�lT2@8w��]����ZtWJ�h<HK�⥞POE `$���^�ٴ�NL@�6����F)�֜��8���67�'Ǭ�VJ��[�Db�ЌR�|�<�����ӹ�,����7��F[#z��;���I<����`�������N
���kjn��z"�AM<(2H��9 յ�f�~㓋�e���wZtg�/�ҫ6ܜO��s��[���?��O�VA�I5��B:��򼴽ssz��d�M��8yt����G�#:��b�/��???���V��k�|��;��no��P`J�=uu��n��"dɣ���X���}�+��X�O6�+U_�}�����$$*ob�	sMq����k3B"��1���]��PW�Z�re��h�F�_ �.�C�`����f��?>����+��������)0��w�=g�.|6%a-��m0�v62	���!dʺ�8�Ā�9�zZ�/��*�ck�d2��҅�?|�J�+b�t�ɥ)L~1]�&����V^^�S��_�6KUz�����_/�	�s��l������u>��7:�9�Q�a:��⩁^>h�ԇ�^�d𗾷�"�o{[����/�m�/(���Z i$��݈�g`�a�ꪣ��J`��ǋ/8��YՕ����6�6�P�>��ݧd�Y��i����ĉ�@Uox��5�sz@���Eb(�3(��N�e:��k�5�}|������� w�D�)K��gd��Y�Xc�����NO
��K��|��ȸ-�=z����c	����-�T�f�w,VY({��6bD\��u��֏����%z�ּ4��ڵb����������<�`z`趯��w&�	 x�!���z�py@��Y�9�T4�wz�2�t�ui��\,nG��E��⫍�~G��~���j�)5�̳S�̄��ϸ����f�߂gO���1R�O�b?��'B�䪁�i^�{{A-�+M�%3dӀ�I���=x���}��xeۭ_����a��_�7��$��cd\�$�r�LCe����@\�\sH��e���ݶ���;q�܃t��5�4G�"���P�jC((`�t��^gN����n���T�A��ȟ�m��ίc��y�ɍ�#d���ji��w����=!o;:"�x�3Po[[�u��J�S�@�n���?=��w��I2v�ı�zF�;�0a'Х'����JJ3u�=��M��>��@Մn�d�P6��v�&mƶ��?�����˹[��>E�IV��_l��]�?��o�M5���hB!%����Gy�j�.�[��s�MN�8"�~��;�n��G�>�!�I-nτnu>�ݵ<�� ���|i�]��~G{�}}}�;- ���n�,]-	�۽u�(�:9�	�ek2��e�=�p�v����#`GF����O0�kB�P�ݙӫ�9�;����B,ڧ���+[�k�K_K�T�¯B�Y�0���M�c,ޛ���ZA1k����Tv��#��~��aPe�r�0�u�_ۛz;����5o���}����& �k�����Ǉm?�΍���i1�1WU�=PĖ�RP4�m ׍B/E��N���d�zU) �6�7��J	�O��z��~,$���ݗ�&��r�O��C0w�-�N�~��аKA��ݛ;���=O���s](�l&x�vk-22���S�o!tqf˻f���� �.��Q$��uu68��$��"Z�I8�H�}"�M k7�n�8 �Ȍ����	�A7y?|�4՝�d�H�ts�c���M?a)�T���� ����]0�?�N���C ��D��C#s��h�z��9�����S�q\4z)DN�<������ez�q]�l]�i �*���__$NJI���V�MaB4����ؘ?8�L�x]r����ɚJ��1��Z�gI]c_�8���v�{Fed�R�"���Ԍ�2QW�3f���8�����а�yrF�|����I����yYHy�y�A��+��;�Nn���}q�ps��&	������7J����L�~<�/r�b��U�Qss�Ǯ�T��S҈��:w鐣_�b;"Z�<1Ֆ�+I����J	}�_B�onK�l`މ��H�����ye�*%�>y��h�O�'K�'��]<���iexj>'hvY�n�h�<u�'@дw��K�0^CC��~����>�S�?�/WUU�w��-��{�N��,�� �T�����Љ�����/���d� F�2.�}�qnƞ�܁"�u6��a[ޯszS�d����:����`�x7��z�0
����^Ͳ�9�����@��v#�\HD|�@��vs{;� �	�kqqqv' �&_dd��;��Ufi����n0O��[܏�>~�ذ����d��.M�0J��o2O��d�*����_5J5�[̢�Ǫ� �+M���ݻ�U�u���J��&�>�Xizv��g;vJ�3�8nݪ�b�($D��J�yZG{�T�8�z�y�-��?��QLw�.A�쪲�%�0����4�\�9*U;��b
���"��B�њ�b�A�q��^��Z�G_74��$�jKL��R�71��M
8��B�� ��Y�M��������F=���괅��1��i�dj�뺻S�D�Km��Z�Q�\Q��đ\đ
�Z����\�}�3�`R]|���>�Y���h:v-������F<b�R�n��}���gX6
�~����;HA-|���Tm�?c�qh�R��
������W^������E@�I]Y�˛g��9���UU���_�ih�T+��uT�Z����O��,,��i�A�=d���Ƃ��o��{��j��� yz�}����D�"Wc |0��
��������������w8��������3+/�F�.Բ��zS��s���#J��%#Cf��"����Wm*��y�v���3A�.ǹ8�5���貆�)�X��ܱɰ�rۿ�|HT�Q�M����
��������!���MX�k, ^y�M�/�L�����`l�\����v�E��.{Ab�k>_��/���0����%>�Bݤ��uv������"/�
 �FԀ:y�#G��v'A���"����s?�}���Q��*Wc��u�YN�WK���R����xQQa���d2�ځl&�T&��P�<�k�{9��򧒅#�|���k���Pκ�2L}`p��0��B= (�P����Z������M����*9��-�ƵQ�
>�k����MQf�ܱ����u��d��'i����iw�`��J���b3W����iAa��.cy#�UJ��5�^��P���x�˴�H [��KXBDE�ތ�<�J�$d�ݧKmFj�N e����,�A�('�������_)�<	��!U���w����~nKe$�����Yc X�h%���7iO�U�E�%��-W|��r�.���#�`I�#y����g~�{{Cg��ꥱ)P�}�.B�c׀whh*Ѣ��z�)%��?r�0�ڲ#�'*@����)����0�
��p��E�p�ף�����ax�(��P�1�NA�aU��)̸o�����׺��h}|}[^�:w�����d��[��2�M�:#/�+Sѳ�4�d��=׸���:ć�C�5$����gO�&>R�]E���e=���[��f���8x�a����P�3
=�E��G�ȑ-S�5��hR�7��ӝAQ䫟H"�M�I��7��\�G��z�nPQ�ç�d�i&z�mc/�3>&rK�ӲE����y��X>����)ӄts���D��u�sH�߯-������v�8� �:W���W�.��j�ta�K�oe���0 �  o)'1Y�fFV5_�s�?�y����og5�u������!!=M.���9H���'���l�eݎ��<k���U�3�	3��\�����w�$B�Te��c9N��~|Zsi:!0p����9)����N��x{��2�ǫ�����_��d��! � )B���@���/������3�Q�V�m��q�!a��5QkiM8 3�\_��ˁ���"�LM#x�c��==3���.&��|���(|����]g��r�9�]��Z7�
�S���/�6a�N�Τ��LO���1r��.�\�%�z��L��fl ��wl,F��5]�>3x�M��rWUM
�%y��Sg�W�����d�O��:���	c���E@q�T�in���K��&�~��?~��k (�Om%��sˊ'�^b��u�	��{	,��?IvL�G+���pn�������a:V�����K�<��5��.�X1����Kj�s��]���󚚙�f�+^? #C;ό������?�z���L�����J���2���͒����E~v<*Q) !�	�#�h����utX=�֟p��iuˡ5@ii�G�>>	H$�EZ��Ť�Ěm4K㪓ӛM�5�m��ý=q��}�l����T�������o��v�Bv:��Na�P�:�xŴ�[u�;���3W�EP�_����pJ��~�9��X�Fw"��藍a�Ǭ���&�Ĥ�����%�?'�Tֶ�ce��I��^ON��{�av{[�����'���5�Ӯ�ڒz���	$��h=��M͍p����������2����ne��]�vr�ů�Z�v�~�,��w?����q�*'D�K`�mm�̸�si�YL[��ͽJ���̻#<BN����`	�
?Wpf��D��|P~��N�a"��-��n�V@'��5��[7!��ϳڝ������4���J{f@� �ـ.D���j�&g��n����&VU��,�F�g��ݴ����0.�r�xH"\rm��[m�d�y�a�G�����C-��q���ݑ��7���YXx�.{X�źZ|X�wq��E�#_�n������/�_G�����U�ۀ�~`�(��.��蜎���1Κ��4���x*�T�:]Ġ6������<�,k�kq���$��P�l	q��OB�e�|JnFh儓��k���4{���VJv||\��mk�3@����WV�A�?ceZZ��m�ԎCk���B���W�]O=@Y���t�1>)��uHt�R�_b,z�.�L�C|�r)�����9����gɄz*���8y�x�W;V�P/G@X8y�~��c��rJ�<?������2��n7���d;c�2)�H����@|.�W	��#��\�۾�t�4�D�:ĕ���;m��}�a�b܏�Ird�%SQȘ�1r��(8���Iw)0!�P\�9���e궡�5*��9''#ּi._u��z�y��P6�~HDY��\Dv��3s�_�Y]M�4M��
;�?�P�V���M	F�]�*��g�խ^��1׶��5A�������8Ug���I�ŷM5浳;8�b�|5I��~�?��Sp;�c��_���^j��K�F�Ts<�6|�܌Zd�v^����o��3���:�n�e� ���HЋ��"I_ 9'g"%k`�{p \|.��r�Z:�g8�Vˈ���ρ4�=�Z�Q�/$>>9�b��v�]�	N�02�	H��������,g!�1�� ��\�%�i �T�ù���^M��SS#Ħ��#��\���-9��A�2��5ZM#�cE���/����� �Kb�8�69ф��+�nL���GF٨d�? �*ȇ�XC�|ӏ01�GJ������I����b�<3	Pf�����|�--�ͺ}l����N�-��G��VU�
������F��+&��ԙr뙶����s�*
���3q��Pc,;�NcQ����㖧�5�Hd����M-��k�����Tb�kMo����i�	�i)s=Z��:�]W�ެ�e�C#����k��Ϲ9B������+"��E�Tо7�y規U�ZFOO��A^U��:Uu���(��<N���MR��`����_��¬��?!_�~�lV���n�����1�����؅�X�s����L�?���+�7E��O����?�GN��7g5�X%BSq#Z�����p�o��Hn琋$F���|B�;
i��2��qNG��:x���!v�.�ʤJJ׀.��Q<%ԛ��E�x|�|��N�H�%��Ӧ���%EH��T���Ta11 S�7�Ą�n�X>}z�ڰ�����+���>�3N�uMM��ޜ�Ԧ��(o����l����-�}6�a��';����j	P1Z[[�e��70�b�f3g��v��:9҈Ny����?I2]1@�X����L�?���������9K]�gH��Ot����Ψ!@Fn�x"���A?M�����q�f���'Ͻ��|lcC��x�/�������m����)�ay�Ӄ��6��H��/+ �֫�R�IV!rt�m�"�F�
~Se�	���.Tڽ� yI��om�/8�zn�]E��C�����(o*��;k�9;���@>��G8)��hh��w��[V�]�����Q��HUV"�k��`�U�O������iNU"yZ��Q�Dpr���CVIf>;0h5U�V�~g�i��K�K\�}�[3��]����m��i�-c��Eؓ�LQF��f��oQ;����AJ��Aj�|�߿�xN������"ŉ1)�m4(�[Ԓ3��Cx��8H�����
'q��g-�	���OAV��Ul�pE�ab�5�K�,[�48%���و���H==�N$@!S�,\�M	?�~>^?��n�Euiv��?g`@w��~/:�8�+uU��d�V�4��D>u�	�o^F�LM5�7A!!l�X�~��ۮ��Gk����s���# ��P��bY4�����Smp��g��4yU��]Oy*������(f]�{m5����ed����2-����u�z6*N�:�.��t��p^3�Q�n�^�3����.7VS[��{@vS!�45��W��}��,��)����o7 �9�z	��,,ϖ#�����[ҡ]Q��U��_��f��b\@6���*�F&���⒓���Y�#8��H|�}����������˰��/�zQg�'� �b±�ҕ񂢢P��[�ǌ@�f��w�7'ɇ��~�6x,�T�F�&���n�z��<��	 �+f=��5H}7O���y�R���Yuq���ܖ�ְ[pp�Cc���8K*�'ɩ\�/-��tY�q������7Ƈ�>h��s1�ӈ�l"�(H��R|��{�󳡶k�)�3ѕ��-���_i�bƁu	6�o����Ʈ�o�VlUlnݹݰ�������������T7�$}�KS.�;�q����S`4�˒�C-�ZZ[�zzdѺ�OM���g��3�D/y���������@:`��]�޵�����|�������M�?D���x�>|$�;��r(�������M��7���B��	�Ma��Б�����5I���ֻ�l�-E��[�t�-����Io �G+���?���KM���0����r�bx���Ðh���8�OK���JԿ:������^��D��ΑDx=��%�$� ?9��W�E^^���H��,�U�D\]��I���XZL���l���P����<x��EQ���8���v$�5���c˞��G{�D	�Bs�̌��$��t���Cg-:�'�����$�w�������1��(�@<$,��S�4:�H��O��'v�V�=sB/��p���,�p��L� N��#k>@E�h��j���sH޳�wN��D+�R��	A@P�.���Bж�5���?�a���r�hZZ[�a��mTU�荥��3��V���&q���sgr��~��7��\�K�X#33�cV�E{��]c��U�*�b͚�O._:t���@��������}��f��2{h�ÿ���Xk|��<��z�t�ʁ)O�s��EV6*n��<A����W7O�AQ�-�����gc�܌U.�@������/�"t��"�|M�Hq���	t�����;�����U���{%$I�$3\3#��M���2CٲB!d%d�nH>�n�^)ܐ������;���sΧ�_���1������Q���5�!�ӿDI�k��(�<�u�l%{dR�@�k wv��e�,�y�|�Gmln�9K��#���ё?�9��V�G�.J$�;#�����N �U��	 50�x�93oؿ�Y^S��1����O�9������ݜG�P�z�V�CxK����%؞�-����Ѿ�cI��II���'��� �8}t�r��Aj
����p �g�cZ�A�J���봵�',�%"ۏ2���4:6��4�?h�w���!���U��+��:�*|��o�d�~z�|wbU �};$9�t6n��������O�Ngo��N�����E��M�������&�r��d4Wrӯ;)���n	�R�Q(m�;��ڴ�K{�a瑱<�g~�*+,�>!�u�.|���0�b�`��B��C�m�dzd�`j�<��9�om��w3;�xbbW��]f��T����g�i�J|��)�B�L�@��1���8�'ov�l nq�4�g/85�B��Me_�R?�9.���7�i�fp�Ε}���<�mNW���-2�Q?1��n�)��������w�y�� ]m^^^R3�\��H���0���>��`�}u%���ekP�!�R�Ӗx���|��o�$l?a�� ���m"{?
�ݤ.7`���+W�"/�XqՇr
t@�qS�n���,�7z��2�5���*�3�  M���u�G�z=$��g��vg�Hv���c�a� ��O�<���T"22!����ܾ[( �0��g���֯���D.[��ȷ�W��buea ���a.bktG8��ݽ�A�
�@���1jd��6MmJ��{����hpe���dʒN�C���Ы�b�F:ѫዪ9fyvF�Ȭi�ɷ�	 ��֭���Ȝ�)�??�<������uq�u�����m?�^�����G�W$��~�=�v�UM�*�#--e��v�����~�_,Sc����,K{]�E��nD7
u]����;�I2v��%�eNO����� &x|\8�P�vv����I,rqwl���E*?9�6Y�� 0TS��Ҹ<�&S��I�Ɠ 0r�sH�gyJfv���,�e#����;&��X��eȠ7��agdp~�r,1$,�Z�W�߀!��WU�kϬ��:�I�Sn�؂�4����ME�$��Z�|dZ��rK�~wãQ ��$�yZ��������\TX2�.�X�:/���I �8ھ��G��W&�N�:/.5+���v�oo�H�\zK�^J�y��h~B�ϟ?5q�{��dh���K�o���������aQn!U�4B+���_=�+��U=����9����EHkF�*�ٞr��\��KO��1���_ݏ>�SnS �v��\�0J�R��"E*�o?H**x��������?�E5��S��!�M~�#�$;3���g�����L�6� �������ָ�g�8�ƆG'�?��0̦��k�F�7:��i̡OCBdt����U�SX�����N=9
KWu���P�e��m��P΍��%�w��׌����:�~K�LI����g������x��y&Ck�yt�}�0ir��Se�׺��Uޫ�	b,��w�1{�����nJ��k8��J�}�k�gC�5�﫾S��k����H��p�W�[�(�F�������~�� U���!��۪��J�Փ���x�v�c��s�l������Lul�g ���N֌`+ߌ,�;;w��D=ԽLɕ������j#ɦJ���_���m{%,��޺��8�	|b�j�9��^F�l0b����|�y0��H�V"�-]�N=t�t<�� �^�-]�P��T��,Sߥ�kM���F�ǯQ����=�Γ���D�mZ�R�L�z�J�RZ
��/LDq����}*�ぶh�������9���N��m���/@�T�We����"/������@N(����Ҳ���>��l��y��X=���tɓ�x� �'�))���8� �{�G��4��q���l[�A��)y��̾��A�ZW>�XH���EA�$/���R-��X툚�1�����l��l� ������s�f�0�L2��� "�K�4_G�P�;:׌ � ���T�{z/�����n��_��֮=��i5>`5_�{q���g١�Hp���ל�V�76{�����ɞ$yf^9ՌT*�<k)�ci����ǓZ�9M,���^/9���x7�@`C�fc� )ҙmiiɜ�>f�c�e9Q���؂��/	�gh"�����D5�qZ�&7O�q_Oxl-aS��k���f ����oO/��{s���$����� �<�T��mdnęH����BNv	�
�?�����}�j�N�404l�ￒ<��v߼{�	,��R��*��;���1Tw��B��W5��O����c��,�o��u)n�z�:s�F��^�{cN�ڄ�����u�@�F� �2s�K�LW��d���*�9;XI. �*�1��/�W� �m-�<n��%4���H[˦)^5�r�w�ܚ�����(�fg?�M���!N�1�/���v �>���B^����d}&߽�$������6ֲ�u��:5G��� �n�%e\�+�"P�y��vوt��/\-��*�0�6��Izzy}�wwD4�R�%:��RRR�<}A�F��L�g'�y�c��4��Ȝ-�P��q�<>h�
w^�y�_�;_��]Mu�`�����uk�YRz�4�\V�"�������S!�W�2{T��ru:{zȁƎ�Oĸ��wς P�����_���G֢�����'��gs��Ą���	������y>�Oy�>�lV9�aLxc�SG��u��mEE��~�����(t����#c�|7�{��	� �JC�#�����}ԉn�/�JA��DN�����JI4�W(����c��A�OO����ڱ�L�)�'
�ؔ�g�`���jӧ�T5��x,�PW�aLŲXǊ�m4]��uD�9� p��[�٦������Y�l�ҿ�* 4�A^A�:.51m\���T��O�)�V��YZz���z�-�Nك�}���[4X,6��LJj��S�����扷��6;w���83�I)�Ǔ Z�[Qt.rGc9F �輦�HA�J��n���B���/"d��+!JR5����ࠟEȜ�e���)�ˋ������H����#5�m��LL:eY΄�A�zIf��&��2~���������k��*S����CBv�����6�o���A�N���N$ob�Ջ�����������j�'�����s���<d��X��s7���S0�E_2L��^�}��GF����w���u��^�xWT8Hh�L�+�ã�����F�~��D�r\�o�6�t�b�D��٢'�����w+(��|�^�G��~�X$��a{|�G��*ێ�ﶴ[���p�<W�2�D8zE���� ]�a���婀�`��b�>
���*�V�Y\������\�o�r�����x��w����NMq{=g}���#%>ʧGBAAQ{#�V���s�t���ŋ_7L��i;W0��?{n��|䴜(�������2]{{/c�x�*��s���C�/Gy�A����%�Jj��3f�ra�ü3�Cn���V�sTT�Ѩ���4K#�q����l�P��e�e���1��s�F���U��9F��ϻ�xn�\��|@-$�vB5~����}x C�a����b�,,��e��m�KR�(�*���646~X\�!�m�c�䔽l�5gZjc�㫏}�r߻Շ����y��x�O�"�Q��H�'�]�ep�x`�k
9��������������U���y<�4��Ī�1��Ҧ�,�I7&�J ���}+��s�ė���Ռ��4�[�� �v�[���d��9i�̹&ɋ�|��TȻ�s�K���b���R*X���265%��?Kw��ʊ6G m����o烠kD����y7��y�#R�is�o`v�ɼ?�a�a��a�<�I|��L����8��r��)@f �j�'4�%���+�����o@?D5#ǲz�Roƕ.JI�ț̬x������<S�`��D�w���5.�9�z9ǜ.�l���r�8RIpf�B�������������N�����	�~��͸��ѿ��UUc�>_c+�ȴ���;�-
5}���EϷ�4o�WWF��>���<�H�[���uO�I��n8К��h��SBʿh��o�9�v�5h��?>M��/���?�\<�p���/�k���m����d}5C������k�^s!F�$����0+�T�'�}.]�|�E�~q�g�̟���h:�@ٰ�*���5_�(cQ�f���d!Q��8MM+����C��^��E�q��&���5fw�\n	һz{�*�Y9yx�]k}�������zڅ��ׁ�Y�����+%��9q���A:g��e���e��Z�W�a��b隠��E�W~�YK"=A�_� �s)���e���nRbG �[8��)4�]�9 �x׏��F�TR�ޓ�^��QCJ��T_$/��6²			�{x�#m�d�\Q���������U���/�C���]H;�ݩ�##S��*��-�B��>8_߆�=��66���ؼ�j�yyr�K=��ov���9^��9Q��=�_��i����ν)�Du*U��"� CT�U�2E��J(���E��2�ْ9���=�-s�N��b{j��i��H�B�
nn����+f�sK����4װ����#�����-�QQ�߽���e[�ջ���S�k.�����T�enl�tv��Q�� ��:��-��8`~���͜�������y7�������%���A��6��*�=+e�W�0�6�Ry���e��>�>=�8����0��kb���[�QiЖ�Z��6*EF���}����C���PG�;nnoj�&=
V=S.��1�z�Ї��{�ccn��Ky�"��eqӝ��?c���� ��=�8�B�[���i�zԽ�݌vـ�G8\����g/��H��殦�Ȣ�x�.G)��˽��֚���yԁVA�r��el�6K@M]�DĮ��[�8�u���9�Z�����]M�]�2fBY	���Kӕ��nm�9�ėX}�}�:��af3���U���8�2���j�VH;D�zg�1$�I���A���ʥ�OF/��ܢQҡ�@#����i��(�4�M�9^�4H/��Q7[�X]$�!U�n��gLĢ$n��ܹ&ԝ� ��t�jgz�[��ϟ�yIxU�\w���my���^ǶࠐPwnR��[O���_��PPs�̝s��������9�i1"%1g ��P��m*8�#�a���gyKԇ?�:^��;Ҳ�(�i-�(�pK��z�� ��Ksi̓���C�F>aR�����|�P+�O|ӯ��1 y.����j4�hT*.���{B�# $�><��C7;��~�B6��=<2H$wN�>��#�?���J��5:4��G�E
��C��E�� ��I�����4�R)))EI�{��d����\$D�h���������=��=�ǫ��x|sBj1%��ZhmP�"L�G�)��N��./<$��]{��t��C֡T_�>�B���K��Zt��������YH���:�"=犟5�Nh�Z(�����@�{{G�oߦ�@s�Qf���r	��9�
h�z5C����3 )e󍅭��(���σ����c��4�5���k;��X,�V�M�>EH��m��͹n�&D�����G���q��7�ϥP@��AyO��H�h�9֌l-5�)ր`��}���7�;8��2u��RV٩��KbL�=�)!-=9q�\�����p�~�4����e�|(M�k� �e�\,1�>>���Q,����$3B-��}TY��_\��A���ҕ+�[��-w�غ���H k����6J�4����7#*#ceGM�_o_��kv�Q��5NR�R��=�\��a!UK v�����Q6���� S.����{�I�	;qV�*�����*OD7�SB٣�A�M��M�����V��#��7��s�\�_��p�^5d��X�\�Ƹ66$�)���Q��h���ZB�z���z$���A���QFbSW[��d��IͻZ��ݵ5aaaP8�G��_���S���$�����[?9&B�>�o��=����<==���Qዽ�e�]{�t����������:t��L�u�q���#:�����1'��G��>�}�B�j�n�	��� �=�3R����a ������υ�U�n͹K:��d�y6|�u�h-J��R���xb�sm�,��KW|��%�}�*0p�Y��e����@�r��0J����c��}�s�gg���~/�olz���
{�T1t�E�[+g���C_��L�v�V����w/+�˥�h_��������4J��5��*��������w�ZB�<f��;���X��!mTH�>�^�k.���(��������7�7-w�@5��ǿ���#>Rn@���@�H(gB&��"OV��4@�ic������.;i~AW��º$f�>���A.߾�b�����Z�k����NH�G/�H֌�,.���ArK��ؘ|e����> Q�f���>s�o�(j�C�TyW��s�Ld�:a1�S6���R z��￮m�������^H5�%��B����
z���c-��-'�r7;��G�o�Uv��	7�����*�ں:7�lĿᗝ�*l/�-���)�᝴ް	��˷�2��>�zP�|�� �l�	@y�X��}�Gi��KK���"TU��!m�ޥ�p��4ܡ��m�d�{�Id�����Ş1-�!R��~����$9�}-|�:@���a��c�aM!�s�^*]�Wn��Z�R)�����#@O�L��a)�Ť�qx�_�,Ss�Q�zʅx~��`F�؛�n��=U�?���<��E����o�\����y&��Ũ*�
?.���N���������+Fy*���c�y/�Ȧ��Yq�[[�E��Ѫ�÷����U�I��u��P� ����s����ES�����9U�'�M:��.����٤4�zђ��u[+��G��v��� ���fz�Z ���T��@yK_Ň�4YQ�F���]Z�=Bf���~-��op}x�<ћ)SӘ�rp�A$~��x"T?|��43cFP�W)���X��da���7er33��"dܾ[~�ڽ`�>-����f?R6����L�ES?���ݾP�c�oO�����c�㬻$R�5��ܳ!&$DF�;���B���泞��mmr|��bY�AWFK�*(f
�>��=�ҟ��.,��i�Z��)�A<�\�$�$�+A��~�G�(�DA�4�:�J"��k';�@�0��R��TFF7���$���]�"<GW=��;���2�F%^k�M�̻�#|s�<2�$���oi
y*���'��h�H��yb`4C6����b�H�Nii��@n��ܿfQ���}x�A��F��{Ș���T�}�3'KJJ��~! �M�����]<7�B!ޫh"x�� 
aD\\]����r:�y�������<T��=�n���	�S=�Κ�G&��p9��U�u�#���7�brk�*U�#�%���~���X�������X�[�5���|�ds��n��p���t�xr�?,zZ�۳tYۛ'^�ʠ�:/elf�;�D��R�Xy��aN�&&ӿӦ�r�=c|�gq֍��W��'�z�
�o`��D�x���(��GB��J���8��oR�OI��!�82�2��!�k7<����9ɩ'�	]����Ty��z@}�$}^s��k�y��컦��W9��7 ֢v��=  ��[��J:ߩ4�EɎ�(��ۄ ��]	Cs�R*R�Nf5���0����sp�Ё� +{�-�Ħ:s�θchHVe t[�%�[��}J?}DL� 	Fy�-F��4�$RL-��>*�ы��1q���jtRAq#@����ne	���z�,�Y�BiJU�C���p�����1�v�� ����O�Ɛ��~v�f�L���eh������y����s6�ڟ*3�`h﷥Sg��t=U"�*f�.X|���oF5��h��=+1n�s��*_bx�L�C��"�$�Cx�\�b$8i",�	"sd��l''�9c��ûl�!N\��~Gq������8IZ��~�=�m���%�Ɏ�v��=�VW���W��vV��lXqqw�X��W��>|�G19Y(�]J��ec�r"��KH�W��b�P4{��y�Ч��Q.��T��3
E�,i=��'�� � k�E�(�򬌅�<��lA�*º����)�����Q^��Ł�f��e]YFrĞ�|�)��n�43����#3�����uY���%�Y�
&''��peh�L��F�r��ǐ�Ώ���,.CD\".)s��4�3�U�xe������3��	���'!wh-��Z�+�e�h�.�$�\
�@�īv�&��)axg�4��T����O���q}��q�g{/������3e��>��^;;�tE�̛7®�'C-��1ǋ�$�b/æK�v�hѓH��<� ��:�$s�*E�������'��^F�?�a��:l�ӊ���v��z�#�s��q��R�����ݷ�Rl2�����{�	kB��Pc+�|�T�0DɃ�^	Vlo�������b����7��P�'����k�E;�O��{r�o��4G�Z^PS�ݩ�w��o��:O��5Uoj.544�\���I��l���n��HV?��ə3���"�CG�!"&6v{5��^��M)ᶏ�:h	6y�T�C��͆��B��~{�߮����>��k~s�9����ȧI��5��hWuu�X��߿g�G�[�]Y�.t����M�Q��1r�q/���ĺ���׳F��L,zZh � ����9�a@kԉ�y�睏n�v�EEӻˁ!6�v�Dw��!����,^��_�
"O���:�X�]T$!#3%>�҇���)�cP��.�8D����Fˬ�r� �%ؔ�3�!ӓ��R���Gꅖ�Z�<�<���C��4�R���w�������M���\�m���B�^M��r�q��jN�@�����ͷK|à%��7d"�SX���	�?�`��3r��ǖ6��� c��-1-�	,q�>$�2���;�H� �}U�\>5��P,���pF3f~���	���pUk�� �r�x��p�U�u���G׸yKyK	����?Vy����T#�����8�3���i�9W�T;Kvzgg����$���hŷ�q��?Kcw��.��V��͜�E��.6ʷh�!:��`��M*b̔�P��"��2ҩ��pv���a򡜞^` R����������'�w�^�9O��i8x�7w�T��9��{�/=Z睟Fq���>n�����2���=;���ަ��C��g������L�W��|��������(�&?����ɮۓ��T��4���%��n���8��-����E�Va���?�{b,<R��<�]������&T��� il�Hz����[;:�rtVO/7��?D��L�λ��_�[�5�����sx�>O�P;%��n�����v�(O<)�wN��Y�D�|��T�'
�,T��\�G��&)5]>��A�g4+�%N��S�A�٢]�)�'8���Z�΁������wD9cNV�~] � ﲽQB��qj��y+(����	�:�C����}�� i�gC�K+k.�Zh�I.C�V �o���H#e������888��{��E��/zά㮸H��>J��95uĭ��J6���f"���O�������)�S��-:�B��������lP���q�Jf�Sǵ<�y�����O�Vb��z�Id�b�h�A���|
l�>�MX#ˉl���U�(-�xd��/�=��7�.�Ą"ύ����A4H4s����hí�Hv�j%��7�t�������O��{���5�z����` uδ]��;���;0_���&�g�z-����%~�Y��q%����TĖ�ϻ�f��>y��٠�/���z��}ґ��V;�����r̵�����������Q@@�C�"�y��BUTē���_g̱5CK"i`�44tϟ}о��ۻubL�c�pZ��aO�q�B�E��/o"ۓ��Q�9q�Χ!�V�N꘿!��ʊN/�<
#bI���LN�) t3�.���8��Ku@6�5�#C�u"�=}�/��!Js���S��{@z��y�A�K��a���i⯬�!��H5`5dB�zV	��,�_��	2���</���ےC�=��Dx\���c�9+����˾&��m]]�����ѯx-.v�"^���u��f6
~�N$2~6H���~0I���Z���yņ�?�H-,I}�IIdΞ��Ӧ�bO����<�_�/���� �x�ÙF��V6��I��Gয়:\��G�i����tTU�Q�Sj�.OMj~�Pe$!)�j�VBi#�\��vQ,���\��tsg�fcD���)���>�6�`y	�{��h�LT�[]��Őc�f3*>��δ�(�w=��^J��	�u�މ&�X_����s��ǃe-��ς�cd���TB�l-*>�Դljm�ս.Rv�H0�~�y���!w�X��sN׿iaF�d��
%On�N�x�\e����L��|�KW`�*S�a�l�B�г8���Sǿ��c��5�V�IR/�H=O��3t�Q<�������\Xa�������S�-n��\��B�K��IP��m� �&Щ��n�Ik��*�����fV�J\}�����/ڋ~�+@�7��Z���YO��便�����c��<vuuM,$`�1r���T��O7����q�$]S.�NN/�2s���7dd�A|ԀmwƟ��9�zI
8kA���B \j4���e�y|Ȍ���Zc����+a	�\��}>���~�T�������i�D,1��\4'�B/���}�{�����Y-/���u�H��0�Ú/�n�ꨈ�+Av�T^}���BQ����v7���y�����W[i�RI^�Y�:= 򷕫O�i?�G�5�nʠbxi4� �HIz˿���A^�#/+<L��M,tl'<�4���7�Í�!T�1��'??�MTÆ&�����P������b��CflU}�Վȷ쾡G�}��_�`6��Ў)�m�L��dP�l0�땫�����Ӧ9��`"�;�"�֢O��k
+��j0$�<O"��!��S�޾�s�ϖ̴����7}1�����?��NI�7�<&{��W�Ξ���>���d�tl��\�ׅ.\��?��r��Q�ԉ� uP�~vF���fcN���h�j@ �ܧ���0����؉c��n�~�7@��MJ=��t�9opm:'�yXn��SݹS��z��YGW��:���g\y��;�R����	�D\Kq1.��s�$I���S典jl�����%��0� ���n��R��k�w��m�`U�`s�3�	��~�3��ٯ�x���G/���&����vv�/��z�n�0~���m͈��RH���Ej`h�;���,"����R�.y�;�������5�Ҷ6��C	�4Jհ�{�����$(xk�GH*\�l����ec��W�b�����FZ�Jj���ʚYX8E��>�z��x�-2h&^�8Gb4FP��
����.շ�HQ��l�>���"��x�-��a���?G��k!a��*=,�oo�HM�Eu噒��^s��1w�����Inv�}J��꾪:$Y#_�i��|=r`�.�F���!�h�7.9��1�"�߬
�Q�P"�ҡ�_�UF������XGU��W�����uf�/f��?��[^�PzM�H!��އ�O[��Q�go��x�Q��2�T��t��鯤[,�r�$�>,"7���i�,ˁ��(oﯸ�_`�C^�s��WINՌ����#::4a��P���������rW��k�k=%W�qd�����\����WMmC�"r�����:�v����^���2�Ts����GAlQE�k���y�V���3�I���B���3kkt~�Y|�γ�z�1S�Oo��sʾ Zg�C��*��d��������-���M�E�*M���
�_(i�1�W�eukF���}���UK_��y�x�t�)=ނ	9�����e�0�����s#5oب4rl�]�F��p��eo�Y�]�v�%t{��j]�������l`Z.�o���-��7YW�)u�L���\������f������(hPd���Eů�P�8��Z�k��A+�ޞ�[X6s��xK`�Vvt�u�[iX=���;�]��0�u�p�Je�5�R�`�b����oC�cD=6���y��2���;���=��P�u�,7EY��~��x�����U>�o���/�5W�#�7*�k���������U	�awo�T�q�=D�+��7Ǘ�s���=y�|h�ݳ�-ON��)+-��̌�+��;��=bb.t'��ݖ��ܼZ�zQah��E�W�TJк2������Ӡ�@��K��T���ہ����:�={
�Y��17E,�xb��0U��lxg;Ǣ�Gs��QXC�3�{5Q�9�G*+{�H�M����ÖG�G�(���p���
"}�;�ǅ{{�tŞ���c�
����>��9�O����>�^K�+�����E�����nHL�`x@�&ҽ�`mxТ�����K���-�t~˔z��ݨ�w��3�W��]>��y;nu���e^:w����ΉrEZ�u��K�<�9�>	P[��ޛ����|�'ǈ�(��lq�q�2�����O� %>*'V����r�E?��Zv�
A�񴂲OȨ���u�]�7��S��햮�]��]Ѱ9�!D)�y�i#uL�4�C����|o��	�����p��W��ǎ݇G6�Gf��<4�U=�r�)��+&"��O����4;�l�H�D���BĴ���ciW�i���׉
�x����������g�w��ߟ|���E8�y�*��e��b��mQ|���nT�2u�/N-�8��DV/e��AV'���"�\}(He?�0?��U/��h��{{{!���*�_�h��~��? �X�s�����4���!W�����K,��o���dc4����]�o�s��l����mFDs��+����{�p����e�
�������FZ�x�>Ř��V��$Z���0I���Hѕtr��o�-D캦�<O� Wf,<{�l�:���KQ�2����kT:�ݳ�yx;��q���<���v��5�ޗ���=6C9�C��"o�p�Ցa����i/�}��Ἳ��NfO��P�`Zj�@��S��� l��3ٓ�|�i)t�������� Dy$�����|�)������2��	.mB��u���ۙ)t�#=����O�<F��S�64�Vz�+�/]�r�P���pJA���&Z7��G�x\����H��2~��IX�&��Gם�TѧhTI����KR�F$�n{�ܫ��&8h���j��I��H�C҈��a�P����bKs���~���F?ۑ^5���*V��uI�+r���2�K�����n�R���w5}1�O���˛g�a���/o�4z��5H9o�>~=�&���,��Px��� o��2�E�Q��G�nRo�qxyyk�X��p��EZ\�wɊg4�OM�/̎:]�����Jn+މ:��������w�Iꖁ�e�
�_�4�^o�X��n�
����`m����(��2�H&�p/얻��ȺϾܼ'0R W��x�/eV���&������?�f=��۷��aD�VUE(L5������U%�]�+8=9IDI�D<�̂vE	՟3T��)Ar�W�1x�M:z��k��M���1=n��ѱ���|P7+W��ip�����o�Uo~r/�ū"ss���i������w����_�V��m8�-,Ш��L����뚠���'&��+���yΫ��@mz�z���Ąb��ڛ����{�{�����|s�5L^~L�� NZ�f�a��]i�^J�I6NN.��nd(������|d���:� @��o��ze�+��
@Q�������:��!A�����/\�;�M#��I )Ҍ�)E��7�cE��+;��Q'�F��_�9"�m�����J� _D����u�N�E���*?j�����;�W���qJL���♖���ݠ�Τʨ�9`�����tQT������~=l���)�+^0(�&�g�:������̏��e�Q�i��c ��Ҙ�G��� 5�mn9��FY99Qx�~������:��ӛx���xc�֖�Q�Y�B�?��#KKO����)���u���m(�#�R��}/}	ZEW0`yZj��īu�3��6��ܱ�u{?��!5|;�n6x�����vM�v��5������=ы�?.rTs�$�W�c_Ot����)��il���T���]]�^ƾ��"�;�w� ���nD����ؕ�Ţ�kj�aD2K��e�p�U��i;��:���gM���Ź$-��$�Jku�⩺^��3�$1��Bl�?��z���d*$$��^��(���hۢX�*� 6�;g@���s�u-�_�V�2R�Rg|��W����߳MB��I��I��S��ȝ;��)�ߊ�v�L�)@w���E1�wm�I�b¸��͚fW+�t���
Q�Ǐ����)���O$�4��#9�3d���Kg�#z��
{5����G����DPQ�Sh�0�	#��ߵʄ����%�j�D� ���2����s�N�~�`0����$}�.]���U��z���t�[�9m�\$��p�����L,�?UԿ���X�ۂz�;_{U�
�GR��`�k�.{���]q[�!૷���}ۋI��J�N�Y�S!d��v*111��@�%�w��}ԥK���w��R��� f���W�kk�HP[�{��rpU~�����D�����'we�;�z�4�N��F ��g��$�D�@�-�ȁF�*���+�6"W��s�ĄM@t{n\�_|N[�+/.����Dn��H�%��Fw������m�?�ϑ
!n �z_���fN����e|�E��&��#��X�(ص
h�aV����Ǧ\��rb8����8���ъ����0OS���&��!����ܡ���`҇�j/J�؆��>7+I�:�����ss�Oό$ugSFK[���u<H�M����Ύ9-�CJ}�m,Q�,ӡ=��u�+�%D��p��(�_��k�T#w�c��?�b�� �i�3֯������c���y��꾖�>/+��o!������S;;�

�E4�\�|�"s��<�c���%�ʅ��J�����:�/����L?WOb2�m�3ر�x���~�mK'�B.�W�������r^[���o�����D���XkÎ�i��ץ;>MOKKc��3-��Q�m�ec���k�����y�k��F7ve��A5Ci�&X%�k-u��H��.iEE���N6�8�UK@��ܰ}m�{$��I~��󼻅��1ᔦ�N��G���Z
�8�<N���P1���/�Z[#.��	��TXݞ\ߙ\��>�V�ks��)����Wo`���J���Dk[ݿs�_^��u��l;I�fH�~u�~����P��}�]���.J���g�J��� ϞR}���'��\a��)�-�<��Oy]��/F|�ȝu�JH����/���tt}79@���Ni��`(;A�;�����V���|����"�O�i?[&�raF�@L$�W��!����h�-�?b_=�q�exD��ۂ���(�F��]�M�[�IE%+M�ڙ��3ݢx���X���\<�y��<�FĂ����W���y�Ju4��}E�_�9��i�c�ַ}�"��%�,�H���ʝ��e�̹�|�c��^�Z���Ž�IT�\;2E����w�D��ӳ��"�X����!
�	W����T�B�`@0�~J�YG� t���Q{~
'.�&Ǚ��r��w]]]��7�s����_"]�z	/zץ�$[0V��9؉�L��n�~��ѣwp���]Ԭ.�}��=�]T �$$>�\������*�|>�#��`�x���)��ڱ��ص��BLV�����d]i������Ab��臃��XIM� ��h������3֞�gdM/]�ߗ���С4�vF6������q\V��mU{�'��������I�'��t��3�7�cPZ؉0��N�c��#e�&Dp\]/h����� ��5��:�g~^�%�m�N���'��R cᑟ���m\��A��,����+��Ñ[$��CDi,�ߥ9���x7<�	�`z�+(����_��,ͧY�t��������w��.Pdɲ�lr�NM�$��pwo0��u��{��A�&���Ib�-��AY�-�	�p���v�~�f���Jm|���xE�C�3����g@t'#H����Av�8�At�.�7u����<Q����^T#t�Xms���0��u����u���v����*nv�&:%�raEZ���XX"��=�42��8z]A�rԳ��^��Z�gh�[|�.p��_��֍̒���y��#�!�����.o{�n����S�Jr�1�<8hFl-0'ӻ+%!&�}��e�g���:�$ȩ��ܾbm8Ψ�j�h��r�EE#����=��"���,"&v�� ���O��{=A�R�ib?��_�H��YA�����{�1v;o�G�Ȇ���I��e������f�{y��;�op�f���2���� �B6�^�s�~ّ��7��<e�����)-�	9���W�V�TBT�p�2���M��%�����nu�x��}@hη���>�����rn�}C�2xl�(���P���?t�r���pM�I��a0�	�)�w~���ș�r*��I	�+�RS.��G�%�Ƚ��c����_�x`�X��;��4䮫<mW<�5�[|�h��F:Eѝ������/j��
[��O,w��H	��*%vv��6j�s�S{uC؆�Y�<S�ck��f�y�~�5|���Φ�<��^�3S��>xŮ\�-/���+�Qr6��/\���a����`8vM6�siI�@�k�M:����&�鰥�%?�p������8�[qY��r[�Vg��x��'�U��ʫ����m�;�-6-� OZ9��:D!�
\o�ȢӶF���3�;/��g�J��Cdx^�8J���"WzO�UfP�m^C����[[��(�5����s�d"��G5� %��(��R|���ff�k ��j���<�H�u�xOvw��a4�X(�GT��_@ɛ7C�ẂIo�֩��J{�^g=l2Ev}�Rz��t��)~~T�P���t��]̌	߉�U��"O�W�l�;(�|��WO/(�u5�s���s2�P�V2�7e1�X��1�{�+��%<2��!]<7.���fy�	&���QdG�h����˛�"�����s�\�	�����;`j�N*0�ȃ׸t�^�ڎG�1#�/�=�+�cs!(rS���3����yDY��ڬ�"8&������S�j�Ґ<�;<Lb,�R�cTYZ
D�⇶6+3s���wl�pT�ֳw���q,��IVK V��.�ۻ���18;�?\j-���m�dvfIɩ��$ǈ��rs}HYF(8R��1(w�'*1!b�NW�����<��-!���}�(�FӋ��!����"B�g�H6��1����=�0(�XN9��9GxԐ���nU�Rd�ϩ���J���(,��b	]�CFA�)���� �m�����!"|�J���I?�A��0�	�H4o��-=r��Ŀ5GF���!F&
�"�範w�x�P����Ҿ��\�|>�Pط_�fz�7��5ց��[����%N{�'�u��}�x՘�c�z�S�]0�{��G�TBQ����ɭ>d��t�1̾Ѻ�a��)�@YTdi5�Tڵ��~|"��0ӶL"k��Tǵں:e�$?����O ,����zx,����RBe'�HI��PJv�ΖU��3��
!{e\��I2.�2B�&�����|����qw��q����|�q�gˁ�\s���3ˮ"��ñ�/�w\�WN=4�[�w���R<��'�Ali�-q��4L����3����|6����w@TN���9?��� ܌����y0>dN�����F��&���FZR�j��j�`YV�f��;��F�N#K���f͆ƞ�ж���r|��m��^��_��2X��C��/,�X��z.���=q�k���^��� �voHepӷ��3�x�ȃ�PLg ��Q,�P���Ґ�vp�L,IbO��~qdL,�KS��&�J��}��e�A٣:LE^���9�M Q_����m��
5�?x��="�#d��BYp=�+Z�`4���PUZ���v�A4���!�Ǉ��>��cR�jV�{2ȫz���?�T�K�d󹗭2w��i�m.���z>{���K�P#�=4o���c��?~-`��y▴x��%-���������U�pk׺QP���b\�4�4�̓�At��nq�$�>�͕�f �i��&�`j������!b|@��N��F h!�$�.U^^�`���[C���!k8�l���%'�O��[�΋a�m���m���Ӿ"oem����76���W�F#x�F\=_�����w����t���;w�u&��/���v�K�w[T��e31E���E���j�|.*J���-J_�y��I��T�)5������EZUu�O-id[_�j)�U�3�N|}|�l�o����qV�:55uNSK��er+s
��j:5^w����ъ�H(�;����� ���Z�K���|�P-0=��HNª�ȍu�z���5��G˩Y�þ�ö���>�y��A�UY�����J,L��!R���E�ww)���l�������MK%u�F�!򞨻i�����JDee����ʜ��`�N{[1H�'���������n�5��[��0�ڃ4��Kn���=y�����6��>�	!!�@u�����i�����t/�3o�s�}�8Y��<{�J(�%��Ը�*7Z��[]9���\��~	D199�S��	Q�y���R��v!S��U*�9�
�ZR|�'Z�WV��T5�3Bڅ�b(�op�BCK+��r�P�ZUٝ�D"QRZ���W܈JW�1��rN�QdM�!��pCs�-�"�����$���dX��"TZ����B����������K-��e�@��2U�8�REȗ�j���q�w��ՠx�&�@�Խ���%��W>��^���.��q�W"�����S-ky))uuyEEC//�荏��ے��<uby��+�HZ� ���8�|�SP�0��~94T��f��=�<O��{�m����	Uh��J�G�Q2��)(��3Y�er~%�ć̜�;��"�Y���:F�~��[.N�W~���r�nٶ$d����pF������Y~&|����|>>�s7�̧�q�*.��$	�K0특gm���u9���?M;d(�6�u
0_C��eSE����}6�o7얦L�
�x��iS��
��@SWiJ�����\v��^��sp<�N���U���j�?�P~��ia��+O��-��25�����&�yq�U��\&�B	S<m��^����[6�B(MN*m���]8����F�tӃ�����K2�$��������c�g�$^��*�ѧ� �xmz���̪)���sN����ww�L��]��DDD�5�\WTf�F����cU��p);��$�p@p�����N�y��h!a��ؘ�	��VWC��h�=���h /��.p���1��:���
��^��ӎ�vT����4�?ͥK6ږ4w}�AF(9ٞ#���'���������k<"���J��쑗�ކ��a�ݙ�;�� ������S���l�va����s���_��U�kb��˵M���|��t�+'v=̵-���8�M�\�)���I;'�o��>-�a�J{eZ�����)i�2'��}d%���}����I��Hq�X�ֳw@w�.M��$s�t��Ȋ����QQ��$'add�g&'���O�Mk�f�T���{YR�W�5wF�-@���TqqqāV�7T+�I�_o�y G봺#������$��'�sJ�T��a�F��-P�w#GG|4��>)�Is��^�11~�����1ί2�)\���ʊ�Ҥ��?���V6n:��(7���<dg/�{���'o�%��5�!��Tʻ|Zr�6��앹>�� .	��+���L�}��z���7X<l��8�%%B ]V������~%�lX��C����Ńmg7~�,���kHE_�xꜝ:p�}_�uO�C���$��_"{5��	1����ȷ|o�^ ����"����T����Ez		��R��|�����^��an�]:)�H���l�3r�we�{m�����Q�VB����nq��A��m*���|/{zh�;��j���C4���'^^'pUL*f��nz�9F����Ĭ3ŝЖɦ�=����555� r&%��.�J{��+�Tc3t\�*�ML�,jci��,�c�{�3�\�o��ɮ�q}�fWÌ�����g�e$㘽F�=���va �w+�����ݼ���l�Z�т��?�W'�[��8�WT1�!�Ȱ����`��d�9����nk�׊���C{���OC��`���L��ߐϒI1ʂ���Rk풙�N����v��z�e��zz4�y�苈����~W++�Ț�Kڲ<�	�]��Y$���5
.ęV���*8�3�߱lu�k&?-idH�'Z�ᄺ�5�����;����ыp�"΂��}vj�7�ODw����~���iE�lZ^I�	���3)K��ic'�5mkI.��ܶ=�)�=�g"���v}=���я>�vN��K߀͵4����B#L*,=�B��R&��R���ǋ�~���Y�_��,���[W�h�u^��Cd����0�QX	P�.Jq�?��F�%����t\�����������L`�]f-��T��l4Eh+���)��cS��Nlmo���|	i�P0���܌���Z�C�༕�O���wR��`���X"�e5)f�e�_ߚ�_��M�	)+;Gt�Ѹ�6g���X��pUƫ7������eh�/�dO@Q4�$�U�@`,�0�g�{�Ė�(u��߿V��b�DZq<Ԉ*p��Ar���8E�����Ld���g|��տ�o:L�SR�R�?9mh����y��ѳ4�ŵ
�X��5�����������É���(���I9���c�gY��}�*��*B:�8��\Ƨ���H�F���!i�̺�Rb���P�|`�a9�
��DK�2�簢��%K4%*��A	��L&��hå􋗵T���6��qC�� � ,�L�
��J������+�}|RL�1���R�������� �k&���Ȉ���mP�ᛢ�F�*�h� 	�~G���5<�o�zƓyh*2���+n6%�(�v��Os"�:����{ɼ=���k����&����wn�@�O�E@�����3F�vF~$Qz��Y�C��u���4a0�_>q$E�E��##�^bʿ[�fp��j���uo9�a�����~*yy��<69�V���!�m�\��ː�N�r��)�cp�
�2硺���a�H􋱅�0�b	��3Ǉ�,�c�ojQ�_a���UP`Y�8������$f?}ͣ�ܿo��[�%����%�>3c^k쟻�
$�0a5q���e��.i�N�f�Ezp�B�|��	�]r�O�=:�$?57S2E/C�rq�B{>G�B�����e wIEE@]�a4�rU����kK�m|��DғQ���-��U�B���>�h��K�։�E��P��''f�IO��FB8%дϘ����Al�M8%��v��X�3��׃�������-���*�gs��/��%��5LL���p��p��T$���ߗQYdi2��:4tb�2눣�H=$��MW"0�����i5�X�,��ȶ�:��M�_J
���R櫙6�5#o��K뱄w:���G�������)��኏��yn}�k-ųW��3���W{�Ï6_K� |�����Y4&ni:<�,�"ě�5���j�@9U�g�O�S��S� �ύ��E�����Jd]�G��ѝ���>��k �fg�(�Wf����;�YJ��U���1S�Ǝ�b}��)�����)���]��X�P�;��T��B<���Tʏ��������6q� ��q_�3�'w����"���������6��"o��V�3���O������s���ع��𞖍�9M�<a�������&�"	�-���|��������H3�G2.����-��<�И񆔪�)�����-�m���x���y�mN$�gς:%�e��p�/Ҝ�Rcޫ�b��u:&������¸�ۧ
پ#�b�l��--�	<D6x��.E^(((�Pp�pc}��J���o����L�N~_����e�<�?0���;#�Z7OO�p#F��8'�$>�������M��A-~���uH����{�Pc����.&PE��9�����`ck+�:,���hd�YpQ�A��5p����&#M�������V!e_���YV����r�C		:�p��d���K i�093OS[�y�����B�̵=�Ĝ+�����*~6Zŋ����W�/e��y���)��t¥�qN�j!H�"|��r�DW�E�Eed�t)��4��I�8S$RY�M�-��&��B#�Y���:n�I�����;YP{1��zD+?���%F�9�pڱ�i"�<���@RjT gW�~��c:�{V�%��?�2v�U�+wŘmf��o������n�{,K�WW�<"C��ea�gf]��07/��8��j� p�&p��vYv�B�z�"��ee����f)U��^�8+�}�`}}����`}��S���n�"&Z%�#������rװ��J��݈{M�]�����}9�ސ'��E�7[׏P/Wʞ����9h�d����2uOh���,שHk''Wfe��rM�GGmm/lz��_�=�{�-i�TR�i"At;3e�EEnU����_5�KQ���w�;��_J�zQפ��MO
C,�k�Ȃ<���m��_&+r7<�Yc���^~':8/�M� A�o߹���� ��UfrR���d�$��q�l`��HZv��U�Z�8FO�hp$��u�c0�պ6ض�翋���"�F�̲R|���Fl������!�pr�c�:���5�Wȉ�����*�yuD��_��1GV�tum���j^��X����O�gCv���kR�lF�^<{��(�s� ���������zv��6)�� ;��6p��xa����l�O^JJJ�V��D�a���;���`�y.�������i�Mtܫ��Nf�������)>�vj�܊G=�� )0Αw��UU��&&�ߌTES)T��+!�C�����*-��jT��#�<L�*���)�Hez��� �<å���p�������N�R�g�E6�W�<HrrǟXXk �X*+�f���Rm���R���u/�2��tI��+�=�� �6����|a�&�71�+�!��KM?�����=��xz�u6���'1����tƏ׋�/Ʌn�Fp�.F�������C�D���%%ꁕ�e���ihh^��o�Պ{(|������ERXz&y�W_�"�����������%)�x9��Kr�QPϨ�i�3�扅�Ɋ�����5�ɯ�(��~��$INGNp^H��#&!���}��i6����DF..���g�(��S<'~wZ�����<���7O����4���+,�������T���3�&t@kt��.����1��M�M�N{����7�$δ�J�N�x��85?�.А��SKs�_����"��of��QSS��HX3k!��+$h���4�_o�ޏk<����<�3���<�	�R���!F^^�ف�4*h���m
��:�.�DHJ��%$������?Ń�D �c�^YAe�̵��&�4���r���5�E!Z�m��)�e����n���aLk����Y��[�3��ӧK(=6K�������kP�/����L~R���V�&���-�sr�*�0�k��t��N���(D]o��P&򛚺
z��I	^��r>��I�`3~�C�c0Nը���*��f�+}/�\�
��Y쑻���HAZ�3����j�BӃ3��(X�+<�gi!�z��Ċl�Q���u�ѥa����Su�JO��+J�#��m�r�8��j���� ґ]�Z��R�����������'�x#�]^�+��69>0 �IOjlmݲ%a���(�96&�cn�;M1�,{f++�%'���B���:_K�p^SV�3H/|�u|���xŞ�N��V�y��M���[L�L��Q�y4�EE���s���cb��y�6:�;�����}|��?p0s����X�&�J����=�lj�N�۷�9[�~�
而,���L�0��[�Bݼ>fO�&�<��J�V.���Y>�n��	/�=�r�)s���:�Oc#��oss<з��6Ų�N���fv����kA|��ڨ�ff����­������C��xD���M��jt���8_���P��nz )���?��w�ɓ:'ffhw�OQ"��>������,H��3���'�,P���,�g�cۦ>���=T�rt0�{���,@���iʐPă�\�JII���M���"���E}$�dʧT7��"���b�s��|E��g��D�C�k$n�9���a��S˘&�����)�7٤�Y����{{�)\��o%Ì���R���=ill�����\��6	�C��	�q�rDF2�-(%m��[Ȁb�=ST\�Z~�n��Y�%!a(�Zy�B���R����;	u6z��n��@��X9$�n2�����^�z�(R��3�*mx��(��\��?ҙ�oXm#8c�Z�l*�	Z9���f/�H�B߇���q��ȭ �����L��
B�R �J�L��ՠ2��ui����ћ��<���������z�:��I���٨#-�t�0��{-vB��/�B_�v\��'o�_���O������F�*�P��%�v�N_	D�� *�l���*�O���/����9�5�4Zt��;�{�VR�,��lZ\�`x��x�FQ���s��*�r�O��t\�5)!Ư�(������<�:�p*����Uف��?t(z�[P��.�O�-���R��`�vBa$n���6͸��v���+/͌������[g�Lx	>��y��FA�����k�����rvKNⶕ�������zI�&AV#w�S�����CK�s��H��",/Y�@#�a���ڃ�s�� ,�Z@X0��>Y ���B�)1Y��"V�;���w K%3�Og����w�_��q7�; =H����1�/8�wY��`z�E��|�J�t��8�=����n�11UG��݇ ��=�����~�0߆c��#�m��uL�z\�q�(��"�P� �olj��0��+)+�J%32��T��(����-V�`j�[卋=��4�.5�Ԥ�tC�Vh�TU݀�{#�|�uйL��e��Op���E��B�c�d��^Bn=�*�`@�����g|��'*6m깭�����> 9Mg"�_@%ي�d`��`�F���3�?������IW��Hj=z҂�D�p!K���
D�\."g��j`@��ޗov�f��~�>��T���%��JRg�.�U*��͕K(�?f�9�{b��@z06����M�.��K��O�Ѕ^E·P��A�AZ��4���8w.fe�_e�A�J� 2��Йc�7N]�y�� ���U�<i���nbHP���%��|��C�؊��y�!	�_�F�pM�i�aŭ�w�^(��#�?ۆf�s	$�6�'��A�,��/��-�Q�p�9-(8� #U�e�������oz��=�f��7a�_K_������?QXߐqcm�^M���Io�Z�p/��$��]R�� xV���w����>c�6�AM�5�bi���FE��40��Zx�	).�|0����ܜ:�o�^�_j�=����c������׌�����9
�x�~�
K��{11�̔����g"M���(���Ln�9�Mc�~Kg�<&��Wc����������{)��B����OMx�e-LpuC�8 H�:e}9�|��Y��}� ��!����W��}��P���s�"��+�U�E���
.�K��)����_�6,Z8[����_���U �&��[�5���GVS�o5���/��n���x)���;'g˴C��������o�QxX�e���������,�����b� g^^��	`�I%�~������,�_��sml�d�eO�cض�\n����w!]ݩ.D�~��I�q�:�L4�^��n���H&]^'Z5I�1?R ;���4 ױo��֊�.'Ϭ���G�]���b�{����ͤ[C���n�B>Ͱ��r'�z���G�H0��&+�΢�x���٨_�eC޾=�I�.�磕��]k��|����ܵ���f�-`+߱�X�_++����Ty�M����6ge��lnz0 ���b��Â��=FE!'"��ڤ���<����TŃiPc�,��롕�pʑC�����!3
Z	6��^��Ky���&d�O[G\�s:^{N��a�lY��@�^�"+?Y�*�F�]SF��o��Uy�(�Q�H���o������^M�n�S2,�����w�l�9�n�k���ײ��w�";��ؤ�B���]��5	|Ԋ�G�}���e��.CV!�%�x��#�<���%���b�nP*�d$-;��c�����bg� ��׷�������C������:cp�z�<�����Fl�C������!,*�C�҂�	B;��`��)+�I�_�g<�z�_W58��Ç�k���w��jZ�n氞���<j�����OP�e����E�����h��p��m�$�H��-1~�������n����Ai�r����E��.��ۯ���sd�m���c���������H@^�`�MP���W3�K�:Ս\�S$�S��SPxc��h�
0P�Q�c��;�!òq�ab ���	��h�ar�������>��b�:#)a��p�c����e�,�ۮ�����''��E�(��;&���#�z��:�d%X�
����8�٧�'9ȉ���/Ȟb��]Uf��qQ�SyCHpT���
�Wk�G��u��ō+�!��u�Qnb�/p���#�A{��4���)�������<99��О�(D�-�s,�FR���+�x�����>�A<w�Aĝ]�,+��q&�2(�X�6��-��.^��x���:^43��%ӯ�]��:3C�l\��g��E�[��N�Җ�9;��)�����ÇLADp�mN�e�����%(�y۸cH0,V�h���M[n�բv�a{+��g{���שiii�"r�Oq��_�@���|hll3?�؈���f�����ψ�l9�F��������������/�yT;�t��EE,�����O�-�B^J�Q.> ������gx�3�J�����}����
��.Xw4fiB�bJih=��z�2���h�O���nBa��o4��?�a��Ɏ9�r/�{���/���z�!߀KKE��v��/���ǧ�	�RHT�iƅɃ��wf�Z{��ub]���xO��QZ�Hx���z��m���5���
��vřI��˽σə.R}J�oB�"�O�59����f���x�Y��*�1]�r�HBB��K���*�b}��i��i]e�jӨw�Q�K�^��O#s��w���U�:��yǆFqr���(�G��%��lB����hV'�$j�0!A+<�qUkѬ����嫸���Ĕ�����f����JW��򔒞2,u|||�>}�[���,]N߄�>����d(ѓq�7b��}}=<��95����~���ͽ�Fu�d��ޭ�t{����G_�-<n���̲�?��8�חUe�m:���XUUPX�I�{be$,<���7�3�x7�`�G�2�_�\���B0>
�C���$
%
W|Դ�q|t���VA^���#'�ؿi0��CXD�ҎM����^[�M}�e9mtd���Zr׫�~��[��ܹCKC��{t��UX��ܯ_�Ϟ]4-��&Z|ŀ�$��������@.��4���]�|y�,�ԤG=wk��*>��Ϡc�$--o
���*�^?y��cs����nAX觭�[�����Og��w�ccMk�<g�+��8���XZO�Pf7�F�P�K��4_�i�/ڞF����0��lȷק	��989y�\�$��Z�֭2ڋ�M󲲮Z��pRX�qg���n��[2�������ٳ�j��h5���x�吿677���,�udb����j>�� �7;�Q��N��p��o o�jaaa���IS��6>A�\��H�������HZF⦲_B�:*��N`������)mos�H_��:;����/��1��@����� 2{��˃����.v���I����D����d̠1�Ztt��<�4�	���������)#P�%��
:�J� �BCm.�='�Vx8:�7������ѨD��!n�;KLOkkM���򴆆���\o�e����u_]Aޥ	�0_X��ţ�>S��3M�0��.������P�������z۾V��(��J�O(�D����{�g�x4s�s��b-��g�߳�$zAp��qB����=j{�>�����L��D-��jt��pr��-~�x�r!�38������������Jm�_�n�*�ȘL\�7M�ѯ�(������m�<�e%��0A�fMNR��E�KaW�n���>\���_�H��L�:�B�s(��Pn�Z�I���tQ+��M��柩_�Z�M��t�k����on~aUWi��:kni�*-D"G ʐc�;�ijJ��ۣm�tG����prv9�D8�������?��>EH��V�F��2K���*�f�^ΨsO�wNI�d��J�u��Z|<�;����)hp3�[P���ټ�[衡�	b�=���h�O��iR�^�=�
��	v+mMty�w����ei���g�f����bi����z��oB3`>n�����`�%6�ʍ���@0��d���P>�C�ml���6Qh����v��-�҂�������[)ii7�;f�Gl������_5Sq��m�]�{���%��ޛu�==ʘ�iY�D-	&n�Z넆���?��-��p_������P�[y:
F6L{�*O���sh��`ajǽ�L�v�P>%%E�� �����^����d�~��O+g�����8�郛/�'J0e��݅�?��ƣ;�~7�1�+���}Q�=�C��jt|��k�{�������3с_�<�����͵���'%��[�m3��y�oݔd�ʏh����G*(�ڑ-+s�c��?��t=,��g�:��A�B��ɚ ������^��:�P[��z���Z�v�+;55W�����c&n�LQ�� J��Л���3�$2����Պ�1X,�Ma���W5M˴@���@�6��~*��ө�h�x���D��bʪ�KR�Y���z'��	H��s�M6^����֖��\!{Am|L����������O�蒐�X����_��o���D�gQj�j�� N��M�[�S�c�8�`|��ring��?��ݿ���L5� �53{���M�a���k[_5r|9BQ��E�X9tq񣃃����.Rny��c\�]7�N�Q�gR[�yW�lY�������#P���ng��\���v>�)����+U�f��
Ϟ%d�8�f����޾=0?�����'Կj�LUG�u�������������-�9�c��}$���O��.�v{�!�K��/loG�G�c���
��+�-]\[Z��sPٔ74�ttt0�L���+�ݏ���?^u�hnP�T�,�����B:!�j��R��������
妧�� �]3rMR��|b��[S�a^K�kk�o��&-�������4mu/��SM��u�
e�{�Y�\�A�;�GE"ˬ��VE���Tء�.����< �,a�蛿���7sww>7�����:��|�}t􎶦�0o�ewwwEC��z'B���\�^.I!i��[d�N|��ޞܮWj�7�,Ĩ�9@�����^�6��ֽ��<t[����p�*u���[Y8����_��>7q�"�ry\��1��=F�<���O�b0��yk�g�t����*J��ܤ������>Yl�v�7Gu�����r�1�CV��1˞$���_�W&�3��w�����.]Rzwʧ�����*��Ν�b�s|�Ƿ��L�=9]otO�����?%J;�x4<�ZpY�Ҝ����uGh�ڏ�o��ߛ�
��e���ki�g����8��N�=޹�QZ^���:��~�]/����u��FHHI͝�����@�۾4+��誷����j
G|9�>��t��x�#
�4��d#�9�V���ް;���:�34�xL�6�o``	��U���|�<����f~U�#�Z�̯!chǅ��������݇U��N���e���l�pq�tT 	��j��WA�m.��tu��n~#�l����]����30�|1�N�9��a/`�@�A�g���ٹu���k��;;9��֮��>B�{�vk�t��M���P�S�9�T����eQ�:>O�{ob�UD/�蘒��6�j4+��L����/-+�=3�;h}O8ݛ&0ci�&[�~~nN�w-�	ZYT� ��v]����*D�<K������#�<�JC�mv��ӲoO���z9y���=��oz��-�����mm-}}#�n����R��޿%�Փ�Eu�w\0Ԏ՝b��v�h��f����W�����e,��~�>7��d5�L��8�#p ��D��N��~c��v�����>>`
E`Y��� &��E�UU�vv�C2��H:J��6�+�*�Ch���:�����EE6�</e���h�e��:���������w�3��i_��˙zv�p4�o���v����o~��d��!ꕝ}M+N��륿<�������<@�aw7ak�e�'���X�i.��J�d�'��}��T�Yj�����.k�YC[��z��_<�� ���xl�4��II���ISB�,>z$}���Tέ�'��^Pp
�H�>y9���ޜe�c���]u�dT-*�urO�LOgsrq�(?�/���f����Y"ş߿���p���tvv������x�V��/^������8[.;�![�>Ꚃ���v��"�[.�����\7���̀��uO��2""��-ncG6b���C���,�b��� ½�ի�����F.��B[u�<c�lml�XG����`J�_��I�2�!����݆��[$[��-���w����f�W���[����/���{���D@P���4��~Q]�Ս�'tttFۜ(�|		����uH�FD��9�O�������*��>3��c��oΤ�{�)�q���Tv�KK� m�F��D��2F6�^�g#g��<�=�Q`�*}N0����ښ����z�O�}S��/�VP�od�آd��ַu�{��z�mQ�6�B���Z~2��QM�; X����e?8��zz{u676����M��:��!V�����6 ���?���`�L���W2+�Kl�\l\t[�����`c-��~~Ǩ$�u�A#C�̎W�Y�����nL�j){��&x
���;����E.�mP�k1z�b���4�lԡir�U1cg^�	�l�6s�����������z�uʔ���ط��ֽv�f�I�n߮A�ʋ��z733�?��=�s�{���@
��� ��)����b�HW5g/r|m��t���O����:Eʔ�8���*|W�6HDŞ��������?}q9���&*���C�c}�%�ݷ�&bZ6���s����#����s�0ߜo:wLT����Y�^���2ۘ�2+Pc3�[�)c�}S���l|R�[y>������N�
����m��v����:5࠻���l�N
Ed!k)9�Bv>>E�����ʷ������z�t1������(�!Dun��fB_�w������b�R��ۗ扻���W_�<��N(�յ�?4��=G�V)�M����7'"b��L�3���|*�y{�u�,-E��n-�p��X�������:e����ߝ�FGF�4ٽ�|��^TП�Eu}؊�M���Q���iW�ieH3Z�����Cչ�i�c<�Nnb4??�Az[ |��M~@	� �[������ŧC[3��-χ��G��1::���j�V����nj*k���5�0��11�4GD�]��G��Ć"�Y�%h;��{]}31+����?��������4�i�Bh닻>��nm݋9���ɛ�ϩ�[��f��#�ml��lwhk�\�Q��d��h��Лԡ޻��"oІ�J�{���,������9y{�_����,�l�:��8Hp?��^oqii�1��b`45��@?�S��}�^���	/j��6��p2�����M�+���BU��Y���«S0�;���Hl�1O�Y͵&�Cu�$���
��ؤk����Z�qi;������|h�
7�V
�Ā%@|8ڪ�P`Ѱ�}�ַ�>[�:g��}����ʬuz�6Om����3���K�D���n���N�KIK=}6?d?}svvU���l5�`�I3�>�
�ʚ���/���:,�>�1�t�����B�:�pkfx�=x��iu#�nm���:^��pB�u�0�hbR������sxk��ϝP�B�����υt=S�8�߆�W�WG���Ū������Δ̞|%��J"�T����x���v����.ӭ�QA���[�@ ��c�w_D􍜤��{`��xs?"��k8���\���d�a|�5���s���X��  ��,O�!~��G��M�d=Ī���`S����}�R�m�,Fn�g��x9���SO�)��f>�t��4�ql]�kae����s&�J��0����
Ň7�{�5�7RM���.JK���v?7z%A[Q"b�=�$SU�o��K�?�r�l{���.��H�/���N*���W�F���x?�8#*���8F�&.nl`E�y���뷧��{���Ò��������G�0�-,`�MdJ�i��Qzw�A��aPH�����K�>�/_jI��ha�ﲮf�>���33#�}fB��*��W�÷�o������q�	���;�f�>.��M).���Ǝ�x��0 ����j��a�&�|Mv���>��*��OPK=����c�ӂ~%TV
����G̗��=*�L��Tp�CX���9�ow��O�[��ȚJ�	��z9D]~>pr�����fJL�@&_���1��P�{^�q�(��w_O�J���_�<����&�sa|yj�0�W�Q��a�ٚ����J�?�@�WkiG^r��VXK�ﻶp�h���1��UP��]�S�o<�0l��<�:t,+`S��׍r��Y��`Oԏ��d�6�$�!��sX��iqp5o��Ȑ�]j�v�dis�$`�K�4�t����eͼ�M�qw��侙uo���-bճg��^������p�I"�90H��Ν�tAa ��ը�*�|�IO2�%�ѱ���}0�K�Shl��@?/�����֝e�,F��������{ݍ>:*G��� ����[^4=�P��U���d%z��5��@/TBˠ �����%)L�d��M�lt� =���w�2?�̈&$1VƩRX+,�a��<6E߶{�h�
GG�ӚnN�|�`��`�H�F�(F�����J���o/;9�����a]��7W�#�������JC��W�C��D�����_��%��=f����D�M��>���:F\�r����]� 7�\�v���r���sЫ�;��*�#����y��U�UU���"???�63�lYK˛�c(K�����?|��ԣi扄���=VTU��ؠqw�o��~:�-c��b����6�������!��k+�4�h3�|7�M�C����,����5��l��C���I���J��ɼ�|k�}0�6N%L���i��\����L���P����7���ia���Ðe t�����-�O�(/P�8p�6,�t����[�D)Q}���*��ޤ�3n�>�]]7.E��yg(��ڒ6��uV$�����U:��z��lPx��כ �Q��Հ/���c���O-|�v�4~�݉�a����N�W_��!�ܹ����?v��)�M͂7�Y��1��R�:%�~�S�}˴î-��PK�qW}��B�p��nS:�� �=8���%`yP�{�d�� �vb���X���{Ga���$��d��ՈG2KY����h�Q�ȯ����uQ��؎�0�l�c;L�[>R����=ZM���|�L{�=��յ�����x>���&I���f"�����vgwR��I���曒YV+XVA�Ap�F��SB���G�q�5��z~I���뜺L��À��1G�%000__�3MDOo��-��w{zEEs'>����p,BZ_���3OL{�T3��5%�J��!�����:��E>{y_��`H\G[5�>"Q��h�{��!/�l��w�n��}\�嚱���k8e�Z��Ύ���忥�+�U"���

0��q���zv��(:J#��c?o%"}��[����>�`Et����u=+^�����1_jO��D_O��LF
7~A��}�'��fDDFV��+O;�t͡&�i T�r��LӉ��V�gCv�pՉ3��+�펙u_�^�<��W٭��T�T�J�7qŨ��)_^P�����L����<)׷��M��R�\�������)' ,`�^��&�T�N���B��8�1nK���,ů�Cs!Qp�a�K���Q�6gL 
���VA8��g7}�����Ľ�:�5�bdp��-;*n�ɶ��ib�}o��P�q��|���`����W�*��>2��8�~�E�a�q�+�+�ݣ�_�����7m�w�Y�O����A���I�iy*BuFpxlL��Q{��MV��d䅔�T��Tm8����R&3J-��N���VaD�@WwwEU��2���:{�{��8q˄�~�}� ���G|���^lb%C׬���a=�y��I�++���B$�H������<�g0��R����h���uT�|����FZ��b۷����E�0?V����r�no[$���SH�ˊ�����s6tZ������x�K��>>��='}��

nn7�b�Ġ�����������[
뗉^U���6O�X�cŮP�����Z�_�
�ۜl'��v����7�~�!��:K�I�"�!KsF�7t��..9��=q�G>Պ߿A;]�&u�E�Ҳ�����g�Oy�^���0����zA�t�t�}�����L�?
5��AJZZ�f�%2�� ��j��e�7ݳ��)وL�߆����΄W�=�����8+++�X���`����G+77	d'������)C�?++�����M�,E��~̓�V�.���o`���U��u�^�Q7p���������Q�k浇˾�/e����Xp�	��P *M�M���>��^��[lS�SBO"��	���L��3�O�:aa������:---�	T��~��g�&�9� �'�q�-*Z�y( ��O�o�R-'!%������f��8�c�4����c:>y�A�G�����e�
a"T�!ST��G������A]==s�]S�~p����{{{��" ���2@��;�\`����:vj��ҡ�pq=�ڜ����Bo+?{�c�P���q��9$L.W�Ȝ�g�Y���Wou�������Ւ--��(Ym�e!��,c��F����졲�J�&T���(d�R�&&��3s?��������ݯs���z/׹�G^O���sD���9��E�.�*�O�3\�V��j��Մ���历_�UQ���K���+��V��������ˎ,{���_=��E�/�QTT_YY��Rl�Pﳼ�jv)x?����D1�~�/�W*Y\<���7%����22�~�2����4����'Ѿ
���0�&��9�2�߅���-3M���]z�)�]V{3'�{{꫰��-Y�9��ⶀJ��K�.��R鶰��r�2 T�^��	}���k���� 9>����a�O]ll����A���ꔕy%�����_��[�{���Xp� ,��t�S�2y�-���,��]ua���}�m�����r�b<��B�{��Tx�W�_�q))))��w�}Ꝭ�m`�+W��}9^SS����C�g�����|~{;*+����|����?:%�+vra����T!#&JO��������
H��
�ujW�*]�P��+�Y2�p�.}~^9����73���0�qQ�"��ߔ��|�/E,���'���c���=����A7;�+m�I����"��::��{S��K���k:�(^��+���U��4|��S�@���:�;^7�����p��>qږim�{Ğs�Xj�aƥ����ɫ��I����Kbmdd�Y��`��������hЮ<�oh�������5O������?bt]�,LP����q��k�+�]�2	��rͣ= u�!���ӝ��,i�M������
�v��y�i��޸Z��ձ5�HH��-.$�z�3o	*�E X���.�������Ӄ�怷�#T(�**Y��K��꒢�֙��vZ��� QN�������}��?�޶�6���ގ�Ћw���KAA��ӳ�/��MLL��[���q��2��銊�#C�N���nh��\"��{�fq��1i��;-������͵SE�Q������O�������_^W�"'��[ZjUj�p�MѨ����f��yiiihK�b=$Q��H��
�DM3s�?�72!c���'��2ԗ��@|���OmҸ�066l�5%���f�Bw���e+���5qў|g&= µ5�?XKѡP(��5�o�!�����ymx�p��l$�Ç�FG�8��GG/�$ܸ���V�d�z��ŧ ��b��*�"�Κ;��;Y$r�n�s��#�����z��ŋw��U׉%�u�%z�&|���;32�]3��6�[d��CX#��D$H�۷o���.�+�,����;Z��(P�wv��Z�5���ɯ_� jÂ_�|��5�p�۷m�&Qs�*��<73CJ�=��4�ɨ�S}�߭}!))�� �o�Q�}��1�Sh�o�^�ݽ������Ҿ``o'?�3�a	��?��e��l-v0]���|�Ȧ��@x
N(�!��v�`X������
>![�}=:%���nm}xK��L&������L�=�������	���Nb8����Ƈ���3�Vig��qx������,0�

�CC�0Ň���A����E?C�.�з��|�&s&�����D�=B1��4{��s�LDf9X?:�<�/��h��t��@j�0�,�iei_��終ώ�<���Ó'������M�|��u��09�ap��	Ԣ<��87�����G�\R�UQ]]ޔ�'��hk;�Yk=V��NGG��ԛ�R8�����@�������� �[s�G!�Ү�@F�FrF���!��x��7T���ҩ_� �=L��!z����V��I�^Z2xQPV�>�U8.s�n�ؾ��0�ea��O��+�k��]�|ܺ�r��M�ߥ��Ӱ���w��"�t۸O���M��C�2��
�k���(ͨ:������V��`p�"�_Ł�{�Aw]��vq��}.q��e/�`��,oHw�X�M �f���1v}HU�zWV2�lٲc���	��))�9D�bEE�#5�K}��Ve��Ь_@J���ˬ}n�"-b��vf)R��)5F�W�Ė𻜪�T�t����__Z^���Br�Qi��c�kA�����h��

K>k�R���atj!#�4q��!9ע��J�By,�|�=��x�&
����Ԕ�W��J���J���[��S^GmB���h�]����Ꙓ��{���©���:��~������������쑻��`R�{Ǩ���@��S�ڟ���li���R::n��t`�c�� �Tq����]���&k�Vʘô��ZYY1nsb�h�/�#��`>'k��+"ӿ���o�){[Ў�!<TH�s�����)W\W���n,�ݘW�=�V=H@��S2,��	� �<�L1���AKED�uu�u�����q2)D[V��O/L��t6����EG�J�j����{D�^��KJv�)w�L�0�4j3O޵�*��Y(S�{��;:���ז������6�6�B`��jk�z�vlD}*���#�-
Y�f�=C?@����uk� �\+�L��C4;�U�6`_���65|���!�w
��Q1w8��{(D�b�L�T���[�0LQv�� |�!e��5c6��t�4�5���yy=Q��Hyd�<�߭T^����7���5s��^p��|��D��kW<�:���p��UL��O��~����穽;7�C�D"m�\��J�E����d�ě��~z��L�4�ş�����ǌ�|�߈�SZ��yә ��Tb����@S��]�9�W�Rk��WU/0��4鉠pɕ�G�w�|�j��/��:(0���̚�qg�g��g�m7�a��X�%�5ƵĞ�ޔ�?i��&󨝡Lˏ�y�v�)�@r������5Sy*������<<�?���}�f�/��Z�����ξ.��;�@�?T���n������y
f�/�eW������g�m��K�C�>.++C���С����������ʸ��6%���d�t����P���jo=$�h���=F��X%_��1Q=~&����a�������k�d�`.6U�^d���ݎ�svt<������TESS��ݷX���+`bll���+e<K��ikw@J��\��G�@vddCj�+�Ϡ�g�Ev1�t^�"��j�ݨ.�Շׯ�AG��=MJ�(GT'�����>���s	�		����$n���`�+�3X^^���7\H8^�����,wQ��@�#:W����ݭ�<�;��\^�����ޓYz���J[�K].��B�Đ��/J5�L6i�.7O_����K8���Ŀ>;/"�J-a�A�}�Bz�ϴ����Ctt��W�u����=�A bl��ӂ!�]��@>�U���!A����)������1�}6{LZ:�'�i�a˵Hc/���B@x���g��<�e�W�d�V�}�n����_�E��ߌ�p���FAnL��!?�=1���$:.�#��^�{К[,�}bb�Drr2D<�$�fvv���t��HN��ڝ�||�R2ݻg�� |;6�t��7�fm�XF�쬀�nW������� X�o��c2j^qB=�sq��<Wa����������r��q[*jj�XXtoڙ�^�	G��%�%v�"�������>H�������+���5��MMi�~ yq8��dgg����±b�.jycc!�H|�.�D��{�d]˗P�@
**�4y��s��^f�F����J�v�i�s�U��Ó7Ng.8�SVV�+F`ejzA��%e�0��b�d���-,-�&&�d��/���H���� |,l
{�C����	��wM��?���tO���6E�]��	c����O����V����O$��~k(-z�[÷�e�	�y;��o7uD�[�=b��fV�<�'P�B�Y�Q8��������������ń��/ttt|����.&{��,.���xT�~(�}G��}!�*G�Z;���)*�d7>a��oĕ��E���̻*?��P%G2[� �-ZP1��}t��E�I�A�D�-�Ʌ���#������d�=�aO\�aXX��̔O�^��ȫ���^	����;�NM�*�`�r�n�gd譴&$����)"MAV9Y~�� ��_��"-�����\�<�ڂ�a)hz��)�LFG���SDFN��sDD�ĸ�qEg�V�թ�隁 >}����w��<o<�������z�������6sPt\���$��X�剠=��L��_�jt�>Ä�K�;s�L���d�,lXEʃ���E6��uu����M�#�[�����L }J#^���8�rkhA�ð�N� �z?[�q���

f����5��o�?�:�se�kj�b)O)�I'����$�jӹ����J�[���D-��>)��7�#����t��&?F�ۭ��r�9����W;���q�������,r� �9����skFx��I���/��5,M�
���LO����ֿ�Y������� 9Y٧���)���T [*՛_@@4�!�p��T:rĜڥ�诗�)!?r���VVBo��F uAt v~f���E|�^MZ��3>o2��8	wx�P�腀�]؇^t��$���l��5��8�dť��@||��ܻ�x��w�2����h�����ݳ��J���[�5�z''ol��0K��|t���jˆ���ٌ�ޚ���#;���1�SS��q��ZG�3�**v����nn����̨D:�Y?�ևd����0��\-D��]�#�f��\K����XU%rcC��$.G_Qe��	�_����m}��5^n��E�xo6���G�Ch���z���Գ�M���::;�_<M����7JԬAz�ZAa[jZZ)�D�ڜ;������heȆ�mш�+��C�.��m���fF� �k��'������ͨ��sX�7�5�y���߾��vC���O,�0ͼ��:L��\�q?7�!�H��������6��:��5��J$t��W�ъA���F�r���o�v9�����J$&0n_IU��ř�!�'���LH[�D�XI�|ӦR�Tb�{yUU����jH�e4���*�tJ��qb|�
��WS.n�=59�T���9C+$��� |��a?�`
0 �D$�[u�-�2���P��Ӎ�Oʹ2ܷ�	�korj٥	8�~�bOb�^�����N��j��G��J>�%�����ڇ�w�UgeYC��ޝx:]C{����nU�n,<Y4��'x��llc���,,�@�>!MHެ�����r� ���͑�ԓ����岪�� �@�����n���Z�;I�]td��1��ە��8��i�����埓�Ew���3WH�_?F��)z
�~��������G��
��/xB�u�n̿�w޿m!�W�����)馼/@/���ܕꔚ��A7�+\ve�Z��C$yAډ�cJq;l$��3%*=G73�;��"� �	�jɐ��)�����#��tB�����l��]s?kj�	d� �A�W�N��,`��D�@�E����Vk��p�"���I�7T�WL��?U[��t�����=����'�v=��u�|��>`�9�H+{�z��^G����Js�4Nt�څcF�>�z�x@�3@����h���!y��v�����o ^Ss���QAQq:t�y�y���
��:~nYi.|`&d�E��BC1���J7{{cF7u�8��b�yA$\��G����,�6���Y^F@���<r:���(s	�����5)��,҇������Nn�k����2���V`H!e`�w�И
}7a��1�f�Sp##6VV=�O� ����|��,++nh���c@fQr��T��׮�G��i+�?��{V����i�t]���Jim��ٹ������7�9!~�RߠB6�ÚC��sO>޸��Ѧ���������z�({㶤{k�Xo:�6��7$��ܢ2�A����{O��$��-a9X�BJ��h;R:GwA�0������P3I3�x��rN�;��gf�7]g:A��`r���]J���_2\co�599�d$V�����Oo=_6��p�v�����/I�\޾��ƙo�jPaֳ��M��>pxG���d�\��1;��Х��ߜ�XN��\�066�;l\;XRY�bĹ֪�S���=wA*����W��oE�*3�}����r��4�$50#�o�Ĥ�z�/9 �c^�`Z�	ߙ�zQW�<�����RJII�0E�&���H����V�-z�O��L݀4ٱ6tt�j\����۠rf`�Zh~avP����K�pkg1�D<���~��ZQT���%���gYJ#�ޱ%Ŏ�o�j+rC�.n}��ME6lx���{�S�AV	�]-'�uSN��Oт�F��ԏ�)%d{�6t�a�	v���L%����'��)��C���r㢽�������s�4���KP��2�y��qE8���DF�Ȭ��^���w��?�V@r<P��`�*~c(��N���]�P�Ha���Z��ZG�i���u��l_[	�eb�0�D��c|ㅖ�E����Ś�L�
,�ȹ�Y Ƛ�"����p���q�s�"�g��!��cW���P��d-kC ҿgOk�D���������~~��IZ�Yu,`�v[�,1F������2�6�u�̟Ǖܻ��:��B\�Br��I�G��ϮW:�2�󖽽D8,,�Z�F!���׸n��+�i쁥�-�(Q��� }ĭ�4] �[���z�V�%w�Rː�Z��l\*����kᓱ��g����96�|�%����ŏ6X<�E���l�/�]-+sY��Z>oh�*O[φ���kR������ʪ����=�X32.���+�M��*ͫ�2+ޓΆI�ɤ����L�� Za��W�����f�10�P^�P���s�E�U����ʔ�e~!���a�Ɯ�!���k��9g���̔��5Ct�(��Ҹ ���[Nf��=_��Í�6]Q�"���#UC�huMv%e��(�Q��-���Y�w>*�B����Srs�C͢N^�:�?VfY�g6cX�����=7w����Ϳ��F�
�K���ۂE��rso�������77�k��L��1����L)��]�h��7�C��o�ml�7����O��p���9�fiQb����v�.ګ�`"�h7�}�&�&z����75S��<:�a����>�7[�����|�5Kˍ���Z�m�S>�.2� 5t7ĻU�������\f��K:v�chu\P@�}MC@>���׶��dz�����0�+����+gV	��0�W�mҸC��Nx��]�^�����.��^&�u�Ndۍ��b�8�@t/;*"� B@����i��g�b�=u�w2P�N�Wl�tK�\YQ[���DY'�S�rqp8c�v0 SR��v���&��gx���Rj;=6M��6�`��1#�0�q&j�F�rei4�Ce�C���(����Ak*�̦�Q�_�}��Z��C���6+���bî��%?�h���>+L�ܔO!i��Aw�s T�8��X)���_Dݚ��n��N���3S�!���:�hr�mr^���O2��͘6�,��~�X�y;Gkk5���3V�.Mt����z`�>f`�s���X7)}�^�	�4 =����P��)9T��gJ��U���֞�!�S��t	UCh�e�n*����E&���u���3ƝƋ����E}�a�j
ƶFi�߭�������V�f�Я;7`φ^I������wz�T�o���?�5_<�o��E/G&hΦE���G0�C��ֹ��e`^y�2K��":��q5�����\��:5�n�5�@��1/�wc�rr��_��q6���]+==R���{�ď[n��NMJJN����h�^=��<��2Ǳ������C{��q�}2�m�r-���ʦ���T٫�cHe�m�+w�k�0��#0���7n�)J���3�*���;8�F-"Ħs���r/o����hȭ��.����~N[w<���>a�6��)io��I2*%�C-�#4��w����l��j�@ ���-&{j{޳�[�qnra��bߘ|真��C�J�1�ƛOi!��7���F]\\D�q�W�)us�ҞI��;[��p-z��0�C}�D����IY@�����M疖�����8�2S���r��i��=��8�D }�T�פ U������;ZVV��\��se�:�A`����<�>�M�V$�-������"_*���}B�@Ƭ@�!�vG�$j:ySo�~j��q���ő��+�l��.��HOTe���+ �c�����aG���u�a%��u}����믕�S��B�DE7��I�'��.]
�pJ��A��r��$v��W�SqII�t~����/3@�[8�S |��0\�M��*|�n�J�cY���.�`�ii� �_^~�Xp�ā�5V]�ڰj����uto}�|y��[TjG��TZmm�>��U	,��ELh"aLV.�@29aD~�bX�`�b �]�6��e�:��P��y��ϕ0�@�ܜ��񮾚�ӻ�m�ҧ��{񌾝g76 �p�ڥ.s���;�ZfV�a����lR^^�����b��d�9C0��kj.��RK�K=��i�ZQ�����WKU�.��E��/$��LT��/��~"+�B��Z@/�8��[�JKKKM}K��㓟�^5���9�^�m���O����v���U��S폱G��ۻ��sF]S���4�4ݹ�.�Q(F2Zt��Op�%)�Xi��kf[й�v�E	�@�Rף�����ܫ�Y�C�=�u�N�1�
�K�4�AG.4-'�!�zN�88��?�dK�~Jȇ\\�Q�o��`���3>|�&n�����s"CxLsi�Do���`��E'ｉ�}�d;���|����	���J;�'�!*QG�l��������Հ���Fy�S;�uܧm� Ϙ�u�4��= R&��{�%�WF����&)ɫ������e韸��S�v��U���ң��. ��<��3p�x��5] �\�|�6��D�iiy�؅�mQ��wv��u�$��qT�K��A�q�%���?��y���08G�(SwZ믤����!@|���b1T�;?P3N��K��9��1��S܊C�xMmu�����
��q,J�5J��6��Ӛ��q��;q7�hGSN�r��&\��'���4��^&1ݵظ�v�y67#��r&�{�P�m����ڔ7u�u����l1Ցv�����C�.������1~�/�:$�*<�FY��d��k����g�v���>|���,V��<G���7�5& i�j��8�-�}��ݘ�Bc_����iŝ,������ݗT�}�0$����^<�Z�x �8Chp�0(Ez�9�,�h+�ZLzH,�fo���Z���;WVyP�����v`��#���R ��VK6]���w�0��u.�q���� 	oC`�{�f�$!������<���twOO"D��l'Q���c,��!��`[a�9�.���:�1ݘy�dB����&$���RrM7G\>�-��]�g���}��f�����x^�S�X�*���=lڷ�������d���ʚ�/$`BL� ��>��J��,1+>_av��l��זa�'S�?9 "�q�\�`�fk�A�z�Y��,/
�1��q��;�����UU/�	
���h<��4����6W�A�'|��]�D��`�7R�b��&h����x�L[n���g���j���]}�"�����*@7�����>���4��:�Jd7��n������
ћkl�젛z�Tk���i!۶�����K���;�x�U
��M�$����7.%��(J�C\�i�Fu�����c��%���܍nd�d��-���d�[�G�Ú�HOc�Ʉ1�R�>��jm�ҴB�	���Xp"�ԧ�Wt��r��Ҧ�A�����E=�E����9�d��������r|���$/���ri\0iH��{;��o������C4��<�Ǹ(gf�\����2��w��V�Q��
khr�6n� @J���k`���r'AX�@��I�9?�O�YZz)R|�w���Gx)Xt�'������(�$��E^�%"���[�U��9��[t+��F33c�:U�[潉}���ht϶5o�M�clB��4��_Z���}����kB�oO���O�-|�p�����y��l�{���}��@�6_�5rP�w"�5���99cl:֛���~Ϙo^�.o�T|�}J}R9-����g�R��G�:yԨ3M�XE^���s*��ey���l��s�M�=P�2(�/f�8H��ĭ�%��	0^� ����:���;��ew��˩����&��5�8h\��6#W������VC����La%�kgJn�+}hb��D���C332�<�'�~i�)��c�*e��(��=��X�^p�m��q�۱���5�� H+���>
W��V�O�������N&��}m�0|������4d��n`C�1����Ae.���q�2s:=�$ȭ�o�B�3�!r��3�w�A�,-R��Mpe��=�o�9���3ss���'�85ni�a
l�2��K�d��h�({[t����Ύ���E�@���^W�1�5������
�Y�by��rG;W��+$= �ܢ�XƩ��y�YX�x��죀zL&��U��͗_p����?�щ󀇰��q�\��<���������sv_h�t��>���,lP�q�D�S��8$���+���N��>x�;��A�AW{�]s��e����T���d��J�ߡ9��:�q�
�v|�����ƻ�A��S����6��Yw�:�ͦ���^  ڊ
|q�����׏291q�Ҏ����637'uJΊ�L}����F��ٿG�CW;� ��
�gE��P�V(���Wң���v@���	fffIN��كt!PV&���y{�-����2��`�
�3!��4z���!t%�r쟋IŶ2�5m�k˵�3�d~Y����yW�h������ҟ�h��F�sC3o�V��d4��5=�\�%Zsgٙ6���<O7|^��$�\�\F�(�d������d��Ø��O���~�T���}�f����Fx�};�����nP�D�@�M!v��s���/�kγ.��q�;��E�!��4��4�.�(���w9��'�Pҝ����#�s��<�:PL\�H,�A��L�o!��)ߺ�X��1����'g$�6�����M�g�%�wSb�'�~�V��o��
�u8�����lsj}�����G&�=��<A��-7G��`�ڗg(l^��.� .yqCa+}�y��q{�ν��ۿ-3$t�������A݌ǀ �V�;�K�ݭ~P�#��b~����w��_��,/��qQ�b�M2������<Ig^�Zp�`��lN2KZ�n�[�¤wf][��9��ZO��x�B=Qx�����q'��΀�hH���	P�Y����(�����Z-K������������;�*w%��TZ��m�u]�P��-�R��4�����i�����չc�k�ux~|]z�p�9p��۰����II���~y�����x#�5�e�v��qp#' �ε�*��`=<,\ȿu�2h�L'^���<um�^⋧� z���;b(�\��Xb(���?������S~�oqG�kٟ���:�+�˕�h�4��t�!�gȜ:�JYWCײ7�c��!t����D�8��uj���N�� �v���n�7�H�*;�U�0�� )ɮu�t�8	�_eG�bz%���S����㲣�N��|�B�b5e�ŏ�0���r�; jb����n��ә��Fe��
DY+6�ymϜ��	9���f�q`sD�I�u��AjzzO*�ȏG�`?~�����h���,J\P�Q4ں?�b;��&k	 kq��e�Ly,�Er���_	\��2)s�o2�����������_K�#�9�#�K���p���S���j$�<�y�:|�*���9KP��� �h���vU��׮ᓚkC�Q�?���J t������1�W.r]�^i�!B��oD$�ġC�\��Ls�T�n��U�e���� ��fN��E�V^�j�D��~�5V���&�����oZM4c����+A��>��)*Y����Ό&��0�X�V# A��|w�3�%@��Ж37��Iڂ�3o�֞�����y��Y�k�-�ί�P}rle�3O5|	����u���9끭,J� 8}}u���9G��(4.��!Ϥe�(7����?���J��Z��芠����:{����0�A`7�؉��B�Vu���H�Ufe��հ\��24s�;�xv�j�������o�)M�� \��]e.D�Y���,�Nf�iiğ?on����s:;��Ԕ�+�ڿ��x��������]��S�//�s���rϟ]�$��ӕ�����rU���	�4�ي�G��--��X��be����z�w�����o�fΧc�J��@�x /�$v:R�
�-l^��Ҡ{�b"v�!3�����o�����mm=��$6lW-YU*�Lh��ts�� �5`(�8㤩9��Z���@�}��� 
�Ʒ�A��!���wa�-�4�WwG�����]��g�7�Vڟgi�����!������!3C�!�ˡM]sb�^;�o17f�m���(�5Ue��V����V�n.�v@޼>�!}U�J�[Tw����G�Ywh�����4GF$yB�V����C9�aa� ���X�ΑN�^k���F��+�L+]��-���<���T��F�.�h ��|��>ey��1�ԑ#;���5U�3-K��cϵHߒރ��A���Y�'���++-�H�C���3M�C��ۏ̪�qO�����
a����m�7^݁Ef"SYE�y�B�O��i��ο/�X��5�?��c�wÚ�-58�Z�B��E�t��`Q�
�vʗ���N��fo�\{����ǆb�! $���D1��,�.r@a��A��d�|�zUI�[�Z����^����1���[�{�K�5�������]���A0=����f�W��J�3�I��ip�-�]�.���d�RZ�R��j���FQ��k���u��ČP��T%K����z��\�DS�h�-�ٛk1??w��Ѵۊ�>��AyT*���M����S�����<5N��e6�y�w��ø��'OF�+�^��b?
�K�I9}}�I���=��/H�w���a�Af�"A���JlWzcB�1�D5�|�0m���(c�gc��
�]��.̟�����Sc�ĳJ���F�)tE��5����|m_�z�k�.Ձ�#{.�zVVZ}����2)Z�M:��؆�'��|)/��[sdRY���9H�U�h��uX��\�B�(�s֫=r^�@�Hs���0����_��α5퍤->��/4��){���s��c���x��C��Z�#4����Z��'��)�*��sd4�]� M �ǋ��X?"��'5p��.�������.�[$퇒ILw��X��U���Z�\�\W���0^�J�_<"�D�fr3ƾ,�̢�����]����� �{ᅬjӣ������������11)~�)���v[d�S@��|�pXj,������V�6��Ufwth��C�N���N�����U98(#���a���6^6t%��c�&
��$wvv�&/�i��>8��ЛkJ��&{�f  ���n������Ǭ�h�����ކF��Y	�Rf0e5�^���J=�����Hk�ng\r������my�M�'����B_"���B���J�⇗/Q�i�p�Z,�FC����Ds� M�U�C��0��$�������VW?��R7��W����Ӄ����M;c� �%��i�5�m��ݞ������p������a����Ԇ�����@�y#~<n;��񀌡��b�R?���M��I��8ŸS�l�J�cP�]ӓ��(k����[ɹ���^�@}�~��L�<2��.�%v[��ac�+���s�ݺm��D]G�J7��ס��C�bMJ��^�2�	��������5�e�����d\�y���(=?$"�g�9Y9��TD����}<_���W��r�J3I�j�ݭ��A�'''W��i��{�T�UMi��*G�`��n�����4�Y������ik�	��._

���u@�������m��\~NMi�����d��<q��tq�f��A�jN��n�uJ�z����� ��O�����7N
Ƞ�Zs�x�~;WsI��yq�����>�)��r���������v%	�ր*	\����M���֞�Y�Q==��"}	��r�'3���J�nd�4}�jC��q��0<�f"�D�A���m\��rǿD��� 99vv2)g�H�rg�$�Ҷ>ał�`q��z�P�Y?�+(tO:-�⣭�&مď�y3I��d#�D�c-�^)������l+Ã��}�ωce��vn����]�o�����t�����n]T!��Ҹh�9��kg�~��6~V M~���N�[<���c�0�����h��e�����(u3�(��������������([�ͨfT���Ie�[������R�m���l����!��n �ԅZ��*�F��!��\ߢ�������g�a.E@CӤ�>S��xJ��Q��nk�5�"��]z*��QQ�wƶ���V����?ɸ�q�6��u��[�P��8} Q<��Hգyx�;������j7F�Fe�#G� H�
�v�~"���J���Ξ��
�>�����f\5N�;�0�Q��V��W�{�A���Y�BY}�\��ˢ�����g�y�W�ä$c�NP��Dp���[�0�̏��ԋ%��"�
�7`��ϲa՛Z�Qsr2
9��p��P�A���;(�9�h7��[���~�n�Z�1�]���^av�_P���X��/�6T��.4srw�\�;B�3'�3@���y`��- U{z���ڭ�뎁PI�y�)����\P��c��3��RJ��J�g�^$!�D�ؓ�iugD>~���dT$*Ǥ�+�5���=���b<�qnrtTz�Fߺo-6cg�����10A�R�U\"5 �k
>�/���p�����$�M��\{�p�am����P!���/�xoo�}̷T���
�5`$�L����7��C�w�2D�ls��)��Vq#�!!�>
���_jY�{/K�ڙ*6΅	߰z���<�j��61x�Z�㌧֍�ي�Sb��޾��V��d�TԄ���֩M�b�������\��h�.|uǺ�L�κ}u&{�y�����[Ǵ�`C'��PG��c2���2Vӟ��$�ס��}�P��lǙ�q�u�E�c�zn2V����ܱc���IvʁMB�E=>>>�
���:.��q#�a�gM�=֪=�����o�B&t0]Gj��^��0��*�U������/0������!�lSB0D���$�!�
�	��CV/K�U>��r��ZL�st�Io�Q���C��ds@DE���N4���|D�1�5��߆��`���
5۴�<�����k�M-A��Q��A��a��:%E�֮;� Fǹ#�z_<�TrZ�w����e#�>�����l�㲓���7Q(j�zg;����(��7��C�X�	���1�����Nv#�n���7�rF���^��"مn��h��B!�r)�\?���������\�Ʒ[�^C���m]7L�,�Gd������� x����8v�C�9\�k�����	����ǐ�Z����9�碷v��q�l�֣u� �y��Um3�)��b 0��-U�U�4�G���p��ZV�@$�H��� f��Oy�|[�X؃�.=��}�m:������.0{l�.�˥������c���d�36�:�1�-]R���b�Je�`�z܌�`k6��7N�)��^�э�������Oh��� i�:c�Z5: �k�4N[�)�W`0*"c��L��˗*\�4ow`�k�)+�����s���}zB��I����	w�y��|^N��7R��o��,k� ��U�tqq�a2	�Vh\�p������}������m�D|}����R��.^�0��n.nn���v��u��i?S^�8�G<����w�R'�_`:s��a~~����?`eE�<��UD�"�" ��OP|�����69vv͉.�aQ:�蛘\���F�ȃ�2K�S�����%jLd������C�0���s�r&�@f[:+`�w�f�=��;7��9m(��|Tʨ8c�W�x�~.�4�s�[� 7�~���>���?|Bt*.�8�U��' ���/7�
�㕠��7J̋�ኚ��A80̥�	�:�②,��4�[Xs��<3�~7���>W��B� ͝;�t��88-����+�p\�e#�g�B��Aki�F��㘃=s�7�QbQ	i������Dͱ�y�[ֳ�8�At���KF�K�Ҳ�=r$[���M���~��k<�F��1*q�2��c�n��ݳ uԙ�[��w�:�`g�I[Gg�'��%X�(�O��W�i���M-ޝ� �Xt�W��K�����WP]܄�c@x �#qפ<�����]W�p�Q���cF!@���5�.| @"Q�T.ϘY].-��X�'�,q���1�5�T�]�anF�;��_�f��Q�Qz&)�w&n����&��kzl��[�8��w෕3M������3���06�ç��f�K�b�B�B���P|�N���Rƅ��۝
`��v������ �=�	��:��j|c��߃.,^e�OP|����Y�&��M�S�!�.��H�B� ��>sB�ݎ�(m�?}c�%D�M��B/?K�5�}B�(2+΅�;�|j`�~x�qqٝ���u��!�f@��e�/���þp�;@�g0�-���4��/�[\�#4��x)�XѨ�؀�~�|�q)bz���ʹJ~����Sx�u�-ҟ�Y0]u��KK��\{y!Hbb茰����Ў̡�!�I��n(���#���B����'��`�:J�ŚW��}�0���9���#Gv�%��s�?A	/<$������qvsS��&�r��o�f`�T=�L�?s��0�1x�b��~�Z`%�������hJ�K)��v��5]����u?��(@��.?�,ݽ���!P,�Δ\Ђ�7��@'2��SÇz
����	T�� �~�����[�\��k��'���X,�?Q�"Y�L8�7 �p���Vp�LD3��f��>9<�9�;��4W��#�L)�Qƕ��1�j��-�k���4s��#���L�2�����֌"*c#
�q#�$X�Qy��q�0;
��55�M\�,��q�����M��L�������;{5�D1����ʨ�	���H$�!�TNO��X�2�����oYZ`YJ��E�k���qS,Q�x�tB��=...�bX�vZ�)�%	Bo-hƑ��ҫ]^t�gU��k��\�/���A���HT��\��\qu�Z���a>�J��I�.p牡X�ҕ�ݔ��o9�RYyq�ѷ�k�H@�_&A�+H�$�eV
-,r�;�"�i0Op����� .�����s,K� :�f;�E�<��II�PNٕ��I��WĆc!@kڒ}.��=^�8��y<�x��Q]�\�E��dŏ>[�/n$_�;���b���K�z��z���Gd=d�_3�&�
�eR�>�@������`�ް'��?���B�Ƭ�2�X�����ፆ>ˌ�����յj��u��kԧ�

�¨4��q��	��^���p$�r��<���~�J�!���r��IT�ރ���OF;�ŸЌ�b�*������Nˤ��d.I+��c���U/��f�3�2s	�ڨ�Ь���"�8ϛ����{��@~M�֩+r`� 3BQjFR�Ad+�0����2��`�?R�=�-���V� "X,777:����GT�7�x���h�,�p�ϕ|�quA/K�P�.�Ԣ���QQ:�_���K�&]�|��n�W����=X���$�1�ƘC��Ы�F�p�y�� �.��E��9fm����B����yfI�b�U0,Z$�=_OT,S�10�,�p} �_=gUE48�Mx�~�Pnn6\V_<ѫ3����P�v�p���G�C��!!F��S8�@/�CȰ��-�NT��zL���1�`fON���$������XA��_8d������u	���y��f�9�]#S��v���_e�!ͼ���0��N�8u y��w�j��CѸ��r>�D|�E%&�}zFy&]A��Ȳt���K�ܸ�`x��K_��2p�jlKKH�s7��ǻ���^9[���cm(└�aP:��C��E�.��Z[�����������j�����&�P�o��t:'�ꤨ,�RT
5!kG!Ր4��![�]�%ˉP�J��,�ݠ��11֡���`01��~����_�N�>��<�}_�u]�������ۗ�((8�δw,4=�.��=��$�\|y{g�e����a�O���0c{�%�x�,F�Ըs$��E���R�l��W�Q����r��������O-��|�����zi��\�ḟϟZ�{A�˵J�.���ik������s���@E�n@gS�t�`t�@!X� ����Ǜ�C�y��⪗[�)�feC�-S�j܏홥.}=5�D�rd�:�͛����_7�;R�)���%u��Ⱦ�~����pW����R�"�<sl�`{:�M�����WV<O7 r+�vt;�̨p�|r{AW���V~��SSץe���־P=>,���ޞ�5<-���-OR](�f6-���۷����	�R_�1{�X��7��_nJ5^�>�Ӯ���J��<�3�+������<#�evzl7��@W�69�G���70p:F������e����Z��h�����1����rr�룭ee'�O���SPg�ٯ��

f����������w��XwQWA����|�FK�6�%=���B�F9�Q���{�[�,#�Y]�o@ա ��=~���D�/>���V�����]R"�����$�v�;,~�|�Xh��3t���6��i�'A�fG�g�K������sↂ٪<I�%QI��Q���V<�����Cm�4�\t�� �[��i���R�tH MW�WB���5�C�j��.|ln֌m�.r���8jh$^����ء���ľ}�RS>����S�G�e�L&�������)
�*X�'��w��f��)Hצ���j�������4N�c9�[��xI�!4���b��,L;��u�ķ+�/�?z�YN�۳����pp���VffG�u�Msc[�t1GG��%e=�����a�U�p�&�m�̭Z��õȘP)�:���9))	��?�,[����(�R-���fJ7.q�r��9ʸ��vv����m���1�����^[���Zt}�����pެ
eؚl+(�SW_�~8[�O~�������v�e������Z�~[qu��އ����K3�ns��?�u��b(���Ņ1���hsf雛��,f�v0����g!�j�"�k���###���ή�.��t����IMYy�C�_}s�����a:���	K������ݾ��a�_�md�#ި��Yd�Ht���8��_9���Y�y4m�T�~�&��J��x����(����w�;$�������=���[B�ޟ6����騘��`��zT}��61.�W�CrHV8q.׽��ͷ�\���=�`�-i��9X�dޢ2�A�|!��(A�R���Ɓ��Wx5p���npf�N�pi�:1��?�z��4�[;<�YO���E��Ix��xD`���S�p��kGr��|�2|�x�Kk��77��n�*���5����NjN��P�/�	�<�4&������u_�^��.6��w�[YXD���wvG75e߽���K��^S`ЕV��a_�����z�����l���@ʰ���6-]*<�@�-�y����� �>�6��|�H�R��iK˘��8��	(�2���٬�q5�[�'--���"s*��|���e�Q���[;?_�����G�~�C����P�Z��yʱOK?'c�Ύ�e��4�طhƔ��o���R��Pz�c�$��Q�W�� bup�a���2�C�5Y�)r.���崲��
boedd<c�=�5���7�v�Z�А:&,�Mv,���~HRrr����Ǐ���-NmF���h�[�Q�=���r����Cb`���!�)���4��@�q������RY�
�M�n�%8h�n|�eB��sϘ\�����p�.�f|2�tjV������m/Y)�>��g_������cr���K��_O^{�89��oK3�M��܌��6�t{����T�E�����X��|in8�l-�"k������D�zW�3���
7�#!w�،gg�ڶm۬���{u%kQ���R��y�����Z	�?�lYDӂZ��Eg��H�����^����|]6�hhd��=��T��\_U��Ko�Z[�����w��e֣tg�,��|ƹ4�|�e۞"�����ߠ�V�雖�qȉM� �0�:�N$PW8 ��h�L,��ޕ�{�Ïa��:0�f�!R���Ac���Xܥ�
ڭqNDЇE�gV��F�@�ViQ�W	���0���t5.tuN?�JN��@�XC��Y���^׎��2,]������V3�����d��'IrǏo70�� ���[M�R8�����l��ƺ<L�-�WU��P��)��			��+6s��D�IL�%����;�E�=(&��N���>���dCqS/s�����J�?c��sP����֣T:;������������hY���Ϫ����0���Z1ˢ"##o@�y�єS�{rt˖-��L�SU�]^��8���XUmWvJ$q�Hsw��w����2,�Ѕ3�_�t�a�yF�7��7pc�r}���l�zuXfff�
D{zzt���_8�X\�rNw����Q�|=S�z�� �d�d)>R���5���֜V�����k�S���ựE�J�<��*O`��cTaٳ�P�x%�V<�9?�s�+�[B��P��c�j��$�ÞL�8����2:5�B�l��V��k��Uה:KO��?dv�����`�[	^���E��;37�M|���g��[��p/Ǡ�6�������+պ_��2�s�#��e�G@�rG��a�.�AQz�;�A�,c�˩��=J�o[���=Z�һ�t�@�inn��X�RQ^��0s�<�Pl.-���
�D��ϗ��G^^�ܒ�B�
��7|�S.Ek����ˢ����������I&�)�^��aw�SL�Qi	)��C�Wܥ������j.�	��#��
��a�{��ֲ�5n�w���=5���^ӟr�'ME�\�"8}AJ�Q��=E�gr.Ͼ���7�{Esz�L�˾�	�~�1��|���|�C�A�N���ȗ���zs7O\7fT��MO_f�A��sK�烊�V�����Oɖ<Z>H)��TMQ�H�25L���p�L�� ������ĪP�+~s�`ƫ+�g^vwuE�R�lk��R*�� ��B��w*A�����$�5���.�>��� �v��s���e9i)K�`�ҍR�08k�2�������-�3����TmV)+�B/0�, �Ɖ� ����rn��l�0�Eƪ�I&��!���/��N}?�O�9�L���V�4���)a�2*T��*�Lf�����C>��kв���]̡Ξ�)�㣇ɉħ�q�'M�iqd��xƩ��L�j�Rǧy�������.?��fm�*�F�W��p�,�~Y��,#�J]_�\nt4��֒rPjh]�2��΢l&���1xi�f%�(h��w�GHY�T�>�x����2x�\ӂ�2f����n�5���ӟ�j�/.yr���T"IoY%��T��\lU���k�rD�a�N瞺Ky[����Њ����2G�S��p��[@V���cJ�-�B�-{K܃����"�A��}�`��՗`�"������9��p����|�����ԪR߾��O��b~wѽ2�g�ީϕ�+�y��uW�*rN���jf���ܣf��@7�|h�2�:�m��Յ�*��Xڂ�k���,��#�RO�H<��*�k���9_:F�O�3��)�s*����=kI���*(آ���أx�����W	A�QI>�����L��osCc�즞=ل���3�VG�7��I#�=��;�TD�2���!ђv�����XC����/�L�s �a����\���(����s�jn�w������@b��`]$sr���I�#���6�/<�COZ��X��z�������e��B[�;�@�2G�=K�2�[��K�SaÚ� �~J%���a�c�lq���C���ma) w��5���<��p(3�e����=v@k�"�Ƈ����82$Z�h��	m��e���-[Z�1��L]�H$Yؿ[�(����˟kn2����j\�A�����c���LA�F��m/���'��Ř]����D��s�'m4���z7X3���a���[AnچZNY󷵎�C���y��Է3_
������-b^�=YM����y�:{�!_��b���ӜRN�mW\Y������f`8G���2g�e���=	0����9%�)�O��LHS�T.����fw�ݐ����m����q��-� �GOY�,�ฟ��HV_6�b��N撓���e�Db���@�<v?�����{��i @>"1H�XD���qֱ�̭������C�f���e�\)0�K2���_�4$�I�W�xE��ѹ�)�֛B�ۘ �M�����nT3�͸�����2�K��?����-G4��b�`�SNqUK*w)�v�dh�ق�T���6��C�u����*`#X�DhEn��E5��O���aҞ9kP�Tql���bs!V�v��L��f_�	ij�0�|��d�j����* ��N�����6u� Z�^�U
�ۜ�rg��ԡ�%�'�	�8�Gų�����&���.` K����H.���TR*9�[p��MLMá3�b��R�u��@���$~��N֧�ݽ��a��o;��]4s ����zCS���qw���<���v��_N3c%@_뾸�,�OD��b��<d�%|�Z�):T�v�p��<�߼\��B��>7����j�CP��{��� "q��Gԡ�������O�×b ��_G��Hj禞h<r�b��5W��7jj�3)� YasT�n'���[ ��T�$�7�H�J�`o)[N����2(=:�C��T �o�t�|�_vhµ�m��r�zL�_�It�����2YdL���kC\#&�l��9�lOm�*L����^ ��dr��@�6��nr�I]�a#��TJ�\̣���M�l���kn��v��}�O`?�n4�.Z�C�|�i���+���>th��� =���[���mFSa��m��b�ZEg\������"�*���� �F*�ڷo�$�t���ڛ|��7�d��������<"'7ݩvwQS9/��i�&H���7o>CH3�K笡s�|���Oc�\��ي�x�߈�n��SZ^�G��On;�I$��B�e��{`�}u@��+k����֣z�ia���-_�0�����D��8Gr0,�e�,NB�ի仱�z�1�:�?:::PrZ�*�҇o���;xh5 �Q,)K�c��y$�K��y��α����H �|���;i��=�֎8�<�u�\�>~7��r�:@a��Ī�Lt)<�+�x���~� -<E��� �R������byH�f�}��Y�|�C��I�xQ��Y�J���4�+�,i$����S
K���S�W��oa�⊣�j(�&#騸=���O+�6z�2�wbJJ$�!Ã�:`�� �H`۾�-����хpD	����1+�4�M�N���2O����u��g�`v!�.��).��ۚ,�>�>�`��򱱱�|7�V�$#K Gndr$Q���s7��b�r��x��i]*�Je7]I��E�x�w�I}�Wz�r:15�#)�M]�������13wF��p`=Г��3�i�R2J�1S�¿�Bר����3���B�u����y�o�P5'L⫂"��m���]�,��@]���0����چQȭ��m&�v���!U�!I�f��`%1ϛ�� �E,�wמ�c��WeK7�\{:vba��v �yq;{ج���?�li��c9�u'� ��7B�c�I=���Y�dO��������z��\s���I�Oʻ��?Z�K��(74����k��T�Qn>�}�Br�aXL6C�����|
&�3��s��;3��u�}2P���q":=��v�Q^V��KKK}���,g�H~>�Wu}b{�v�Um
zڷ�	= ���~łf�녮}ŉ�Q�[;L����Id�ʞ&�9?rNe��ɮ��zG ત$�)8�F.�K��R�LAO����3��h�ݦ���#ebH`�����"����8z��K��:���z�G{V&a��	XCG���3ؑ��Z�.�.�4˱�è+��0��M��������v..j���ٓ/K�MU�}S5�[1_���+�W�#����%K�C;OD֘�#���m��0P��]���!��a�D�m��;�`�ı^8�T�¼,B�}=��T䕖����S;�r����

_����\�F�x�� �Db��-�h��ύ�&�/�{*��O'w��+�Qp�+��ܽkT'�!t6�57߆a�?�n�	zMM����)+<��s%��zx���{�0d�=���Ѹ�M�!QM:�+H�Z�����H�=B�l�ɧ���C1��Q3��*�>;Zjll�C��~��JA3�$�U�B�E��o�儭�#Z����x>_��aAg��+��5�<��c###K��T6�
iа�U�b���#����_}���s�OvO��)���>����)��Q��xC����B�PŹ��ԎLIS ���y�>���i��D	�P��/����t���Z�2b u.�mx+���Yl��ɰ����9��C�o{��.��
I��j��kj���<�Z�WQx2%\,�cm��h́���Ka]�jʽ��� 6}A���0�O�ݠ���UZ��[�B��=ox����vQd���� �W"P��h3�9@�%=�T�#����0C>���Ta�|�d��^j�M}�r���Y�9�899a��Ә��F�1�X
��`�,��,08j�e���PV*n	E�5;kh^��� ��U"�j�权�i�f�!;�)����d!TH_P3���<o[D ��r�-�F�FTH6泲��f�� �~�x�)d9h���9i���M-նe�ݓ�0c�9%�C[�b��~z<�9�3$��G����+��J�*��{XB����"<�hg����7��p�֜��yR�2"�,�� �u� |�`��y����j���g$�%LF�����3��T�RUZBf�U���l@^�����?�^2w���$tK]������T��5�������(Rهr��S���f��$�J|s�^�jtv '
º�x=�I���"�Vh���|~llj:�t[���X,�6=V�Óo8)�^8zKN��s�$u*��1�xE�:$�G}�A�nBЏy�ׯ_o6ʵ�ʗ����#������̊1��caX�"K���̈�4���n�=vl�}Kjtfff�A�I֞bW���X4��c�[#r7 \C�V\�,A��XZ�,��Lj��
Z덠��ĭ��{���8:2���y�b&�8�r��_ϣ�t�� C��ya��Q����6|�y�Z��h�ژ�J�j�E�@X!Ơ�<&�~��VӜ|*Vc����V�^� �Q�YN�·cV&O^�P��~�s���IY4�?[؊��h_��v|�'ߍ�,:-�m�oIݐ8ӴY?:�20 ���fC�7��ֆo��+e�`��ڮ'+y)M����T�
����/n�S�x�x��	u�s�E7��+�o�)sH���!�����9tfu~�C�����$x�fc����jV|�ba��M���5����I7��9�4�� s:I���C�S�rH�N�ޖ��o߾��"K}E�\^�>Q$t�v��f���b�(�~-���;]}A+e���0��KE��*r�:��y/�]}J���R�2��6k(����������L���R���v������dȰ���w��[�l��z���R�.E��)���o6,���a9,��7��B$@���S�uN�eW�5Fqq[Щ��W����� #�\�<����^��ȅ_�Nf�*�z&����8j߬�ډO�*Bf )}c���˧T���`�4����XaKٱe�"���J�����8�R���oR������;�p�	��)�mԕ�L|͗����M��������n�p1���-F��s�[w=���([x�5�O'F">>~�s&��B�2���5��F����GPS��AW|��C�&[�Ғ��1�� ��QdmAA:�U35��4�`�Mi�v!�`�m�t:=̙����B�oN�W���A6��5P2��W��7��ʨ�8�J)	�7��qO48I�?T�6�Ec�hcc����G4��XDh�UB'�h+�3��ERw%FW�?# :p��e��
l���VM��;dGd���i\���"�����BM�!��<�ui�4�s5���H茀'p3���j@;��$�_44��y<L���cͻ�I�<ͫ��]zْ� �D:ج��n���P�����<#�V�L��y�V���q��?ʓ��v���]Ͳ x;x��bL:O�4�=��Q��crr�3tS�n߮E��$h�Tx�q��?���ؒ(>�	�HRH/o2�c~��@v�T�4oA���H\'���^	��!�]H����CbKx��4x�si� �N� & ���W��6� Fwz�����ox!�&F�!�BO;�8��: mU��7Qh=Fʖ��H&#�����P�Ԍt������1�W���V�$���|��s(YX���ί"cf*��5t/h7:x���E䅈�16�.#�S���A-̙^J�>���Lf9%�=Üa袣��>�45Q*�(:�g/QW��0q _��M(P[`�1�����
7�hr'�Zy1ncq�}���N�u�OCCZ@�� '9����^�ɕR�Ţ���5��+S�'�ƁS-�4��ҭ�b��9���IJ�7_Ns ��_����.�Bi׉e̡�)֪���f�y�&���^�L�@(�̃�e#[��P�fr��	��"y b�k�f�_��eY����嘬��
�Z�4N%�������M�����m��vq�CZ�7z�,��I ԠS��Lt�-f'qH�*�ů%ڕ��~���UC;��G;�z���9�rj@�rf_8�= �f�G���A�Xc�<𨁽��ކɛ�/l֋��ފ�f�?��&gp�ig+�\9P:1hah�5;�=��a�#"kdFŇ<u6���J���&S�SBvb����/�XRv$%�,��ma����5@O��������\4̥��Kۙ�T3h��9]]o��E!o�d�-���"J�W����8����s��nʽǏK0�@#/��S(mIc��)�=M�7<��;��M���>��mz��P��?JI�RZ=�����h�H�N%7~=e���J]�UR��ۮ�V|Sq�3�T -C]�_s/��`�����o~K��ޮ�d��F�2y��b�*_ϛ@TNp��T|g���t��>0�a��ѶPK4F����O�@�%P˩�u��ϼ�Yӳ��~j��fP�~#h�5O)�A�T���n����i��}�YUt\\,��S��U-6D^���Q�8�9l�'�zQ�����h��0����l�/�a���|��R!�E:w�k�I�$���p���K��ߨ�	^�[����"�^t�O��nQ�:�B�A�!��+A:��)�Q�a��&;Í}���%��Qp�����&�B��;w_Z�0p#�7h���1���[$P?zb�$�X��k��5��e�sO�˥�2�`wQ_;O0������GS(�a<�t=ЍX�ޖ�b��c`e�)
<2�c�s�}�����Хu���o�ai�2Yq3��n�T�k���x_9��ߑ��]�Yn
� ܔtceF��w�=���M�͵��HZ��1�_��"]�V��KA��"P��,�^u����T����p.�*��$�S��St߽O2���K(�| ����u�@�I�����r�ѫS���HA�V��~zQ���C�Gmm�������^}�x-�8'��\�A{���z��۠�pG^���K�7�>|�l|����q�X�k�pE���*7w��5��&���d)�7�P�P��*�P1�M|����Fݘ��XR��j�z��9x�L��H�m�͈��sH�E�֠�"?5A.�r���̲�O^����04����c�S=E�x/p�D"t��vO���)�^�x��?��!څ�����wM$) K�q���ec&�����!��E^5;�����ҫ����?�t��B�o�������]�x�)2%��/64 ���3e|�	���A�����z1ϛ�GC�����##.=��G�����/b\{y�,?�`�\�,ggϰ���@����՗24׶��~K�s3���c�-��Ik�=XU����JMЬ3�B뻌���8��P�v�-w��<��]	�Ç)�Og�^8$�.�t�-�Q(*.��G��-����L�R�(NC���Z{{}9=I�����A;v�D����������s�J�/_�~�����h�J8��)?� ���������@��X'�W{������]��H]��`*�`�w;g���ƌ�/꿬����I��m�蔾������ݻ���-BL-p������X;5u�իW�����6u��F�Tȁ��pHe���
��D�B4��j�p����P�H瞲��ȪJ7���%��_�-/-�$�3E��"�* ̹��\geŶ�2S	t;���`l��7Ͻs�s�:Q5�q��-@��K��X�bYK���9vnmoo m?+˹�9�K�ڍ��bK�� V��s2V!1yD&�c�>�k]�N��5�x���ɬX�R^1�Z�F�������Zu�Q:3�	���^�~��T�nW!ڐ
�\���'�G6˹	��+�Zs3jg~�����[����+�͘܅�n<g61�6ta	��$����ccو�����.SB�p�!����:�ؐG ����h�L�S�W�����ܻwr+�30қ�lش3g��Q�o��H���B�~�7��hȏ@g��gdr�uO����h�kE�Q�+&t/���##�%~l�a�-X��e�*��6 ϰi3�Νhra�N����Wхc�>%wz�3�{�-�D`��jM�A�D��!�=�GBSD�%ٻI
�5��#����U�%��ڧ�*��]��#� I��� �%��Ӽ֧�A&i������Wβ���Y�>6�8�T�wuإ�s��?�l����>�D���ߛ�9��׎<a�Q��M�_����p;����۽��?;�(⢏�,ge�rTC�d�2�� ��*��꛷�p���sO/{~?���?"|��X4z3�ہ�
����m>3����?_�ϊ�yV��ܝ
.W����ꔃ)���:K���!e��Ȱ�Txw��^8̏ѹ�H�� &�<��c��D�B��I�J����Q@@��H)w�������X�EC��Œow��P��!�RjJ98[�n�Δ���П;�a���s�8~�:]��f�I�"�8�NH��ҝvr���BX^���� ֣����
�C�������j�E�tg~�G;ٞ62㐸$�������6H�v#]�82�)#�5Ac����Չꛎ���zE#���`4�"��(�`~��{I3��L�����~�ey.�{������-��7�m�\rڄ<).�G{Z�M�t#�k2�O�������eLUnWK�R]i�����MU�$ü��v��BS�ΝIݝ�S�᷿ߕstu�SpQ	&s2�]�^��s]z2�x�9sje�A��=���Mr�M�IB��M������
�.|�r�K}`+�S	=c��b^{�\����>|J�8tW$�GsP���Fv��z؍�]>�6�ٱ�ŧy1p�S3���K\�'.	�L��+GZ�ǣ�omTA���@�u+4͆�k�?�4Ìv	Y��j�/6 %���-#��|���J�}��V#l��R"����wd��[�{z�tzΔJ�b���
��{+H���c�9������^'�\��ܾ��QϤ,7�aC�]2w�N�';��/>B�Z�E�h_�N�w`Wa��NN+R��������E�'~ExSY���D8�� ���V���3�6ю�I)\�2��UA��?i{����	�m���6�^`��o��In�n��Qx���uQ�:��D����F�k��Đ�נ媓(tSe�'P���t��y/3��ր&@�(�;�_>��/�rrr"֗|��رa�����W�̋��{�tKWBRR�c�O���{n���9����V��PwO�U��;7�;�r^me�����ߏk�/�<��`����$�#|x�tc�u|<g���N��d�MJ�AȞ�	@-GN�����)� �pa�2t�_�^��"��'�,C��r�c��r���P���1UN)����u�^���\]�b?��("��]�hq4�B1���V��)�|V/p1��7�qP��Ι(~/��3��G��&�!frYJ5gn
d�;�6$��#�--U&$G�T���ff�f��K�B�EEF�U�l��~Kkt^�z��"��a�ֳ�i��Җ�4c%�Y.|���3ߧ(����Q�/}2��F;��:�\��
7z)��q�v]���?f���ţm���q��X\?������t��'�Vm��5l79�R��e���M��|z�&z��)��+����>S3/�1�Y�?&��R����gc�����,/X'ly�����f�#`yϮ[v�&��Fi��X�f@>B=��u;"��I�CP�I&s'0*��Qo�:ۙ����:2���^B��@*\��q���O�+���pn�F�W��
q�_��閗���**&f�U��Q����z�ZJ39�K�Ts�\`N�xȹ����b'���I�����LL�@ЪƓ�����2~���H���ZVU�BȎ3x��Hj���p���<C}3�X�E���ˢ��<cI+�K��D��6������i�;���ߚH�Q��ke�u����O8
*xX���	��cޅEEOu3�D�[G@նB3���޾�i�0�6d���
��+UyP�@u�D����'K"�N�O���U�i��	.7@IE�V����O�f�|��Q������!c.��5�1h�Es����$1v���Hl�e${�F�Yvq곲,T��d^*��vU)=镏�o�N�%�V	L�d2��# ��W����Q�τ� �i�>~�W:�����3�1�Q"�2W}���h.��Q:����ë?�%KiM��u/[����-[�Eƞ+�"E0�*W����B%��3Ϯ�KoIN���g(��t����?x���t�N\H$�m�Y8�Zdg5��q�\�^6=�_����XwL�C%Oǜ�s�rsp�Y�b?�8d	=QZx0���)���j8��/�~q�Ι���͢p���(�#k����W�*�Pt��v)��0>��Z�^�r,Bn��=(��=�_Rx����&��_1q
Ӊ	��T7Z��aip*q�t$���rv�0�砂}>�lX�����?.Y-.�H����z�'�B�	���Urhׯ��i�t�A�l�`Gw�?�꯶��I���V��'C*~я�Ȩ����?�qk�>�c���ۓ���l�5�D����������H�j���-��S�5�Y|�|�)�1�/�ʸ���o$���!��l�J�Y�_��M:WEW3���58yV4�X�q��������@4��3`O�`�׀P������� �
:12�-��5�:ѕ����)K]�;�k��!7_�ۤ-��k�˗uLx��U��u�^�;��ļ���d�)9v�=~�0�i��/_2퍝��M���g#x��(��4tc��f�u�F񈴽mD�v�gm�[Q��}��7���`�s�5(�LG89�?5��U��N������acɢ��k�[2]�i��PU�|G؆2"k?�,s\\��/���j)�Y��B���9����P�#U8����G���J7h���#��1 1�n�Ю�H%�Ĥ���!���ѡ7�dj�<p��J�Z;�s�qo��tb���i��_Me�/���e�ݔ�D��������+�h�Q"��T�i"I�IY^��_Ey�:3`��xD���T`NpU�ڑ9�[���̘虱�)T"�#a��k}�[b%�2<���{���`hVX��?|	��-�kO�&S�{�;S���~Vԍ�QMh�BT�̠8�X�g�G7��vVcmFj,i8 L�3p�	{�x~fpvq/n�ߤ�Z�z@HH��K�{���#3� ͏��k�{N�bA��S:mxbq�An1ɻ��)�αTV�.}�xU�*�l;��^�{�	�Z�ݱ�H�|䖛Q��Z��*���;��y�LJ�a|p�X�cEs��L�i�9�Q�֓�>�֚�}F�wtgH�[�!&ּ:s[�s+�_A����n�O	����Pȭ�d�����~��ʅ�OG�;�L��A�ڙ�`���_j|o^T\|Q�6�a��W�H���o�2����ATO!��5rg�)1�/?L��ib���z��k-�9��Kh>�	��&��Q��w���P��#���Yo���W�������RVl����Vh�X-�4���q�+ב��A��N/g-�mpz�5>]9r�>�F��i�M6PSxI����a��y��DED~�E2�s�a��Nc=�~�		<RWٲR3R%>���d���\�MD+ʾ�u2��$j暛�knް+x�%?Y�!1�����6;�q��c���w�T�gDl"
:��9KNMg�+4p.B<ƑiM���ͥ2w��UL��?Q8t#�_����*����6���!�����U�u����z�Դ�y�pAI��ݝb1s��Y{#W�4*�	�zjiXƏ�� l���)��e��az�˯��*8;��$m}XA�0�����*2)�!-�$.eF��q���L-|���wo�h�Y���%��A����&��\�]��í���t>1_���_^�ˍLL�������Pfo���/!&ځ&���D�����(1*��f���ڕЂK�x�U��G��3�q��o�	Pu02�ӗ�B���G����DFOs3s,,342�h���\�P�q;v{t��ه�j����]~HNh�+������^��G��`0��E��G*)��绰8�k�j�o����vI������qP�'�����䐩&D�e���37��By�L��@��ԙB�B{ky�����]��0�"qkB��[/3X�]�-T1����m�**���?�)B�m�l ⫟Q@no'�:��y^���rv�(Y���"���h�o���05�r<A|$ݨ�T����4������2���Y�mA�\z{��D�Aߏ��d���ޮ}����R��n�7U@C��� p��Z<��GF[5'3���k9@���L�R��Wa�������5g�N�����u�۪�6��gƚ�
FNW�&C��|[||l�V���L�np�G.y�V*�d _��Hx�g[ak�p:C��UNь�;!��/vrқ�_ p��8��`%T=�{u.xI�7�͕�͠CSf�V(�*�
�I��;��@~5)�V��ΌWg�Ţ�;"�;6�1�P}����P�3�o�}�^6I�1 �,��p�T�m�޼��Ј��� ψ���͔s{+9
u?Pl��L��8k��&.D���z3Q�w�3���j�3��N���64�scn�������j�Uq@v�U"c.-n�FX����+���}k}$�+�q`�\]�ſ��q��)ux�dT���}�D&�x*��+�w��^"{�����"���$�y1���)�e��|,�5C��l� ��_�{Ї==Y��x[ۈՇ)���z��|���#0F��٨6<P�ۗa��J�-`6�ҭc$BbH�YC�9��VV��o�wc�x,�,������O�9N�G.��m�꜇��G�ޫ|��� ~�� ��]�~�����7���k��������Ti�s�b�E��	��g�����H|h��IM��j��+��#�mޠ^���&��sb��+V��$"�R�uw}�O��X��+wwu�{��+��ۥ�H�~��.�]ۏZ���99�ҍ��s'�t�:�XR�|Bn�H�?(�f{{�����aJ4X��\�m�Y����Y�T�򾧟�֔j@�
é�Y�u®ً�ń������Qr~�����	n��Dl8s
�ܔ�EF���X%�f$����͹W�ޣu �촥Д �r,�P��!���^SKsprhs���9�JV�	���E��/�w��|��o�>�����	ݼ��§͋W�8�$��k>���!�]DJkw����z�a�۫�˦�M>h�?B$��6S8�	�TyV��G	��ߗ*�����J��o�`�zD�5��@���zb(�+φ=�}������G][�T�{�uM��N�@!{�F�׍a��99�����z_�^�g�rή���qx��K;ِ?z��emܥ�yU`hha$891�;�7T������"u�b�Sл4��mV��@/�%tE�[��]Z;B(��^�����_Gw�Ә��������e<��.U?ې[�靀2�ҳ��$m��,��p�o@��q\g,�U�q����l��,�e�]���ЃR���ǯ��?8c�$�Tq�_yU|6b��K���4"&�S<d��s']��9I��{a�mxA��u(��t�3�IVu�Wb�/Mm8c �dw6���/[��A�o�\����1i8$vZ	���T�r�[��j�,h�|Y!ˏ��Mꄡŷ(�N��L6�J��/�T���s*G�Q;@0 @Kj��o%��x@�Yz�	�����}-lu�]b�Ui�[��Gaq�w�H����љ�%�lH8ʶ�OrPJ�p��x	�6�|�:�4��8�!��zkڧJIq�:�r��'TT�q����f�a0��ݏ��8۫{u�lv�2��i/Oz,=�������T���Ф{|�%�z� �j���nVk�cն_��~&�ދ����l��W�[ �)���4�1��V��6��Y��)�k�r���3��-"��|R_����aa~,�7)�	�Ώ��m�I��#��v��I.p�ĉ�]�S@��kmZ!��?g��ӹ���^F��,����]��uRJ*&��(?K/i\�3H�#��M�u�_�EK�ZG�p�HÞ��Ƭ�Lf��s���B8��_x�NH(lSpo��0���o��be�!������Ew��֛fi�O><�\�J(�㶷�z��.��+��8�!Cdu�.��&��ۮ�G%�=�m>6+}4�B��.��R{�C��
�:�$G�/8�dw���&���~a��^���]���\�ȝ�j[�7��Y�O\��@�/f?���lk��m��}�3y1m4�SH�X�Ԡ�ڮ ����MQ�����+.��3��:�A�I�[�W��>�󭤆~���3T]G��Y/\��]�w��^s:����iOq��Ch���^���w��O�4�S:��x�k�~l�?�
T�'4
�>�|�Y��7-�!��q��\�8ipN����Us�m�c&��ܺ ccc�!!zt�;S��na6��-N�7���3(�U��>g�jao��1>�����r!�fuɟ..�U^=�k�/�s����|���G\6�?����W��ЇuC�#R��G|�-	��S.�/�*��Sl,\���1\�d���"&O��>�F>����[�5���ĕ������==���$�;�4�7}K�k�^�P�NP�)�b���$~�n�͐C��}Ƞnۓ��o m��|��jϭ��#k��gf��XK�г���|稤5Xy���'��kg��6�9�E|��*�#�:}�(5���U�YG��W3��+��nޚ�˝�!p���1z��
#��jj" a���S�f$O�̩����$�Z��&B?ޖL�>��6�Ρ1��<��k>�J���E�2h�p�@�1��� ��'���mU.�e�Y�A��ۛ*���J7��$@m���DCcm��>K[]\�q-��p)� Mv��B#�0VCY��j���S�Q��5�lIrv�H�K7�ןݾ�G*'�-~㙣H���\���z�:>�f�Gn,*[-�����z�K�YR�j>U���y0��t̷+Lp���?6o��ٮ�uUQ�܎���MiG�!�1u��ſ%��Vt|�x/��6��ݕ[��,XGE<李EO�E����/���_T�S�'[��������?��b��j��i����꼫]���WK��,�z�tds�O���ѥ%J�y��lՐ��9�I�<�R<��\WG/�8�z������Yͥ��&�EUà]��^'F�����T4��6i`�@�y��NO��w��.�{dš��>���&/�����"
�����o^�cX���;���&6����\IA��q�O}�%�CW��<��O�i�-��t���͐���2��B����;����7��VPGA��ڈ`T�`1"��A�����Ju�t+̈!��!E�AJ$JҤ�B��|?����u��de�˓g�g��>{�s��O�r8C]]ʮ�bRB�깡��ῒxju}	Q�y�v��b8f�������g�����Bj'�'`�ď�4*o�J�z�Y� ��k>����\���w�i�VVT�}m�_�Կ��������N���H���zK��dݘq�?������̄=~^���O&R�@Җ�	�Z���4��5*�m?d��`!�)��<xw����A�Zn9�Wk�rKl\N��ݵ�%s��T�U� �ݒ7O�'�x�Q(R��!~	��6[q��R���~������ ��q��m@�F%b�C��"�>y�x�n�ҫ�tl2��ϙ�� FN���i���,~T��U��e������ߞz����Q�8��E|Ɖ:x8�" �h��:�I4����X�UV?���b��ҡ��X����g�r�������g�M�i"6��6�a��7�G�S>�>Žc�P�w�ι��r�+�/���pE�����C�����+��8شc%�Ĥ�Aȋ��f�M ��S�+_��^�2���KQˇ�"�yp�j��Ɍ�d�({E�ZˇF���-)��C�r~Or���]v��
�+l���FVq�&��\�/�8R�;�Ԍ�p��rB�"�=�_�խ�)KWX���B�N寅t���W ��Rp~�5�(~v�ο�4�X/~�Yu1qI�'�F2��$cd@��)Z�^0h'_e��ysGҖ+�ޢWazf���q�����++��F_,N��#In8�&��}O7H��J��#��=*�ͯ����Љ�2d�������$��~��NP�DR�k/9y������[,&���$+9�K�d�xV���aYWU���7?vA���։��|�`������m��Q�J��(�%�n���Uv�Ck�i���1u��Q&�w��>�(�Y�ē=22��,�y��zE����@�az�
ӗ֌_*�N�#/+��1����=A�?�������)�F�  }�yW`5�����7c����ٸ)�p����X���������ū����7 8���,�����7ъVnٹimSp��*Bȍ��۱�G��J�g�d4w�f��f���(ﴃ��"��@ 9{[���8y��f�/v��tCQG��B���j�Ҋi�	�:�
M��ϰ�q�ħ.�Q��,��e�{��
�J��u?�L{`��-(��*�1)��ҧ\��$+�� �J��Z�5Oe�*5 �)��p�
�.�8{҈�!X�J���8��b�%���P(^��?/�]h!EC���H�UͿ��T���]�@�d����t��?��7�8��BFX�z��)����m\r��� �dL���I0w7����A�HUA�eV4u^-���!��`�Bk� ����U:6.�m ��K B�d�mB���,&�-��A�9^��;���o�1?6����
k��:��_Y(It�!K�&��@�p���d��uÃф��Θ!e��H�	�G��ς�ZQsk�����%�C��N�˻�:$ѳ����
��w��F� �� @�F�R�<N�cF������Q}�,
<��w�@�$��SE��
H�F̃n?����ߚ7�0lp���c���-	��f��,�R���/A>״��������6�����0-�M
<���]��T<L��e}��s��4����俗�� ���a0굍q����u�e����)�+��/�� ��R� �+^��U�����ߥ��
��}_���(`8��e�`� A��t{�P�����f���!"�d$�z��#P�]EV��%�9H�EUz�pӁI3h4Ȓ�f�$jf􏏏?�J�A�b�Q�F�9�uG�\��.��"��H~�։# E���ws,�-����u���w~�	,�����1���l�-埥�}si�-�m�������0�-���A�h�%�P���h��;Y��#5�֣,��\��	`!��~��G!E_>K��O:� ��ew�nGW<�'"�t��Hdu�D�p2o ��F����]�.�� >(I2(��dl��j��Au�wVՈ^�Q�m ��������ʎ�:CZ�,�ͥ���\w�3����� ����9�@/�ZrabtDjU;���8G �{��$¼�4�;w$Q��0�K�oP{>!�!k������	���Q�M_o%Q�뭴�n�+nuY�@���-���Af�VEE�n� �TE"(,N����J��f�UR��;|e��!��bEÚܵ&�$�e���D�~4 ��dF��`��&jNd��1MT�6��:�!g�e�M�Z�f䡽ԅ�~��Wf�s�%KV�^��]��ݘ���+��9�_����ƹ�Y[�;Eod�d�-��e���q!=�	��ȷ���:/|�l����Q�`���D�MV����3��W�#�fe��D�g��S�h�`�N<F26}�yz����G)��dD��[9I�U}��%%%`є�H>�#`߆�VF �2x��൲ׯC�Z���yvDYE��"b���Z1��y3*��]T��n�Jj���qR����ZW��*�b�˪u��M��s�ٷ��6P��F���WA�Zn��1�7+Q��G�Y|���B��iI���Ew8�G<�.>T||n��g�?�>������J���y����H�Y?�˺��i:q5��k5�#ȆF�ז���}_������9�\�!!�0�k����Ю�HO6���g+{خ��F[���猪�#�������{�u��K��������QUo0�A�R��ؑݻw{��@t[��N���s��3�֡��w��2��2Լ\u����p\RtY��[W��F�M� ���nj1�ܔ��w�Fg�v�Ai�~�֚�#��h�)pzF��D��Y�t{�+��k/�j$}�%(Iw�[�~&qX�{�Jl:`�]IlW�ߞ�����@��̈�.?ᅗ��<&�#������>9ɮ!6	K���pT�)@�Ź)�����@��޺×���ȵ9���d�-�qj>ӄ�ϐ̬A ZK�����g��@��?��O�#N��3��neHt����}�K���׏B���$P<ӧ�{����,Ev�m�3a_�}���z��v���98{�w+���Ht���Zc��F�S��P�(@��0jT?Y��x�$M�����I)8��0�H�آ��Z���ĥ��>�X�Q~���ē U|�<��:��G�O����>A�������}�A�}���5��3�^��-�w�<]�bʜ��RZ/+�I���=�/�jż�V�*z$�v�G9��f@Q/]E�!�_9T�:1�[��=�U�g���-�3�M���ǟ�Aj}��G�����>$���?��,e,�L�� s)����$yb$��Z۴'�������"�J+�,w/�lb˩4h<�����4�3?�����A`�Q� ���*���9�\|"����\ 	!����Q�ɸ%op�M�>�X�]�ԛ)ZZ>���6�V�ҩ��[;��1��	�gAY`�h)���ڥ&0�ϣTY����܊
ڲ���]�O?׳�cIgh��s��>�vfa��,��c��yg��"I8��>['��T�~��T�.
�T��8�I��͇e�E��u z�Y��ݐ�ġ�m���|'�
�kbd�A�tz���$X;���_��@�:���;���ӸUrx���"2�:��O>���# y]��{�
�f��\�}DMf|�&~���z,`���u9�����<j:!�5��K���9 �X$�����⑕���?������}�|z�j���\ZÈ�6�$H���g�P�qv���'^N�K�~"A��(�ϑke.;|�����C�#�������d�Ê�! ��.�����~�W�]�d��	:{�[Q_��Z���b��+U�Ϟ.6��.c�
Q��7ܬ�>r�jއ��ˉL}�g��,�7�p��*�ɀ#�[8�xH��}IFyon��M޴+�zk廍w���ξ���_�,J�BK %���섾�`�q���lɆS��YXu^�I�kL��'vd_e�1���GC��Qr&��@���o���̓�a��$&P��L���0���LNN������}V��5c����/��ڋ%�2��6���G��Րj�.x�G�c/�ս�8��0��_��8"񘌚�x��k��6QD�z�qR�����Ꚛ���oQ+�a�:[��40��6��a�>�u}i�}��`�(�\q+1I}8 #��j�NuA^��ێ���݇�?�]w�Դ���֧����Iޟ۸�d;$�2�%?n��Ã�@����;�ۻ�W�f\8�&���k�&T�1@�j�D��c���k�$�O�8�'������	C �H]#���ߍċP���D&��� [gk��m�ȈNa!ǝ�T+����h���^�٢�F���\)_�zw��:O � �jx���<�niI��OL\Zٟk#g��:E@��Ja*$�s���H��2'@�	m�-����%�Di�c.DV�y��L��f,²���X�f2��0����K�Ǐ���2�������ك�+/�?Ǧ�3��*�-H�1�,�-X�(oB��1���0v����u���`��j����kpDxxڅ�Ja��N�W��|.^�s�U��ԙ�I��dm�Z`[�����ط��U��"ӻ���']UrU�ML8��n��7ͧ�����]0��?�V�WGf��g��͝�ԒY�ل�!�����b ��D��L�K���!�n~�C�}�8�l�8�gΎ#d��ޅ# M()+�����˫}���r*nu��p�U ��z��g��Y�Y����Ӌ�)bEe�":�
uk�=$�=�Hd3~��W� ��4��P��GN�ED�NW��7�ǩ�U<	�������#���u�;�Gq�j���l8�^��n���4a�7�;�~k9I���F�h6u�pp�i]��u�y�39lƄ{�H���nؗ��"���ܟ����`�1D~��G��#q�HksI�}]��3PAX�C�ѡ굆4�ӟ1.�)�W���<�i��NN职:�*M�����3��+��.ɍ�9�w/<���S��6�U��"�����u@;}�	/�������	p&��{����]���2���[��G����bP�G���2�{[�����/3����?��ӃhSki�ㅬ�[��ܼ���>�Wk���V�?D:V�u��s���ݸ�� �V��5.�a�q�j����'�p*NL�dG`�9��0D�s#�u׌k��^�_l��Pd��UL�ƛ33a��ᣥ���3���{{��Ig��&/�zEi��]�7k����"�1õl�f7{��O#r<T�rz��ʕ�����0�z*ֶ�*�'�-BM���u�q}�����ټ�0�@�-)�LV|�a����	L�X�s����oe����4[��s����Aov�S#M{b��c����v)���:��0̞y��[\wM�$�5!\���<�QK�b *�2�%�3f��¶�f�z������bj`]�%�E�\$�n�����#�R��n1��� Ѯ���mq��9#��z �<R���V�a"�\�;_�ߔ�-	!]�j��!��ԫ�}���{��'L5��?�1���Ev��VF^8�^�2��+�\a�	C7�ٗl�cT��\Yk���6?B	�2cц|nf��["�
�u�!�c����c��M�%h���OR0����2�hJn���]sA*�﮹QT9����J�.�rF����o��B�7�n��VDTe��Yԕ�]3	\���	+���CSʠS�����g�p�Z`�k.�&�c&����>��D�s�R�ʹ�U���\x�!|J�Yr���{��"�s]3T[��{W��G��;Iv�n�-�Z0���BVe,�ZA�g��K儚��!L��U��'���l"U�Q�`�$7 /k��m��:\�Q�a\_	c��[�2��,���
��{~sl'	�NĪ|�n�$��"R���R�YفT96y�1��L��c\�O^�f`�a�{t'Zź���w�W=�B�������0"Ùb��W)����NDF:�&�Y9�{j&�8���:��j3i��O��g�h�W��:��R�Y-��T�e�
�j�Y_�5yY6�z�j�����<����h�F��Gp�uj�pMÏ�����ܑ�D�� ��hka�B�l&��b��]L����V���Ϥ`+3{G��]��-{yxhTd
Er����"\\�[��b�z&x�Ӏ��%� �d����׌���6�������P,o��Bp�7����n�ָͤ=i����X�Ǽ��1~(zt�(�SƈL��B��:��6��[�g#Xmq���DI�T��Iʈ^%�Y�}l�cH
 �񳙰�����g;�J�L�-�^"�����Ԏ]ų�=�T\G��wAQe��!O!8�
�S`��������ͷO(W�M0��Rnogg�p��t 6�'$�8w�=6� M 8�ʁ:j�ʪ44����(]F������Ʊy8�q��f�<I�-jD�&Q����俟4iT�|��~���������X*�D��W���N=&�T8��čj����Ij��$�I.�\&�Lr��2�e��$��/�.�C N�f��_&�Lr��2�e��WI
ٍ�N���;�qC�Fn���7��8�j*´��ҏ���T�?�~���������#���	.\&�Lp���gs�%S?�V!���I��<��Ҏ��Do�C�?�]r�r���'�k�Z��&�~4F�+��ѫ=��:��BM�L��4ū�P����$�0�Q��7K�:أ�-��#y����/>_�����rI�:�����j��Uc���e��UI�?U,����;�(��Q�=���÷셛=��D#,l�|a~��� PK   V�X.D��N �M /   images/4f771273-f62d-49a2-b0d2-ce9da7065853.png @@���PNG

   IHDR   �     ;��   sRGB ���    IDATx^Խw�\W�-�n�\��9��j�rN�������`��8�`H3�G00�q 8��s�d[V���S�X9��{k�*���ޟ��>}����u�9����k�V���p]WS�����/�@yP��p��몫VAmjک����e�lջ��ܛO�#�)c b��&Q�����ôl7TȪ��OT��W�@�4tM1G
�,�)���EM�,��uM�#��KJ��)�^R̲������@ST�Q�R��c�m���-��j��+��p�K^?�Hs����{�)JY�hpm�*�KW�r��Wo0Ӏ�e7��>�P}�G3\G��N(l�����z����r����ݏ�z]����\,_���Ǵ
V�)�ڀ�h#�eem�l9e�q��*�b�E�lY*L׆�±Wu]KQ��9TWq۵ǱU�qt�,k����~�q�vt��*\^���P��]�>\> ^Gq��
�[���X ������ .��N� ��؊m:���xT�Qt��g��
_���J?���UE�{�8�⸎��[G3ߧ�P]W�!Ô���
��SWuશ���E�!:.x�2n�Ǡ�Y�w?�[ރ������*.f;pm۶����	�*w�.��#����Y��*28��F���+e���0u�p|���=�-�����^��3_��Uɿ����a-���/B�����r(�J�4t�e��A�ۧ�MN�bk�m[saۜ
6��3丰iG�b�PhT|�P�(ނɝɽ�b8��	��3^y�u.�a�
D�����E�"V|��h�����*�Ů,���{��4yO�}|��︼�7.�������?s��w��
E���~����N�����%�Q����2.�Q�i��h��m��T�J?&�ͻ�^�Wo�\%e�~~Z?��P|*\łj8PT����CWB��\����o}��׆5��o~
��;�.��7 ȕ�t�ꃪ�a96,ג��E��@U`:&���E��tE�|Oٶ��'�����1���H�(�\Յ��Py��*�$nC�+{�q�ٻ�gl�������voBu�Mc\��s��-�7�7�~V4M&�����-Ck���Ò��F��������ާN��͕���υ��gr�C�U��bht9ޭ�������7&~�c���x�P�/�*���*st�r	�h��/����CP]��P���;.���׼�O��O}k��f�:��̯�Wu.�z,�@��`+>�5d�]%���hP\��z7Q� ��F�}�	14��K��lۂiZ0m��ϻ� "���qm86�{����jr�ғ��\`N�<�3,Nn��8qܻ^0���"rs�t1۴��S4U�ŀh�P�IW
�J;n���AϪ����g��/�_ަ�,�L�G�^#�b�/�OxޥjX�����Q����-�獟�#��b�g�jȮ�T�ƬҎt��`:
LK���&l�N� ¿�hA_F1q��7|��\{B����C/�����,�*t����y�v.L@�`�>X0�8>q����딠�TG�ω����W<�q-Yx>��}:��M�V��Kc�?N�eY�B@5Vã,�Fo��İY��i�=�ޡ���cT<�x������d�+!�Cu�b24q'>$�V�j��/�x�=��BvVé,��P(&��r� ��`]9��7:W��*���ÂK��l�дx��p�~hzP<����:J�#Qǲ0�|���X�`+�{�i�n��'>����uq ����x���K�`����d"0��i��AB�N���*�,�0M�E���`B��r��{1ޒ��B�`:�	x����4M�|GTZ��	��z��zᰂ�*����'N�����L�9fU�P�$^�|����W	��=�:f��{S�
�*�E�����M�|��2���{c(�=,'��X���:bpm}���H�M���,�a�%X�#kcZ
J�[@1���D�D(��H!�~+�͙sn���W����Uʺ�j�����ϯ���4\=�-�
El�N|c���+��T��G)=�P@G0�O�ñ�J��V���0|(����kP5��)\	eUU=��jH��Í�tR`B8��<�D�ߋ�d���ǀ�౐s�d3T��D�.��,b+zX�x(��=9^z	I�d�&�@o�Dh��Q�mZ%xJlZ��4f�%�웋N��&|*����F��\��8 �2Ũ�V>'�/���|�F&o��$�X��U�\'�0�P ��!'�{��n��MW��<��㋷���wz��[���n"0`[z\��F̡�
�f���.C��uQ���LR$A(A ������(lYT_6�Z �?�"3&zo ����(��C��7��ty�d�Ъ�Z�9��%4 ���J,T<�Jl��D��ӽI��	r�KU��D�\�D|��@�(�,ج�-Z�*��tPe�fއ�g�C=��a�JV9a5�P�H�*#G	!��e�45?tAJe��hi�Ǣ�31��S��$���t�r���cמغm7�����H"���CF%R�"�i#5�������)����-�_�w�U}��<���~�k��bG����+irc�l�]�_�0�l�P˖.ĢE���5����(�
AO� ֭ߌu����A�Զ#�G:W��B�<�7����.��&�щ��8���S�*���x�ޛ`�JXa�_}����h`qԉ�K���C ��*�^�j��1�|�� ��V0�ê�u�Ұ&�?1�����U�"�>�k"���Y(N>�����1kZ'��N��"TC����ЁT��Ν�e�.���M􏥑55��A�SP��[�P�o@/����n���|����ӿ<~��O����,��b���B���@PC��DmT�E��Ι�\y.����f�2d2){���H�h-
E��������� k�K�PU�P|O���x#ӱ�q,��������D�êz�
h�~�a��&e�t|�ߋ�d�}WV��1��FTI��4�������z�f�����=:E�W��M�K�00.b~E*�@Smz���ҋ�C21�TDMM
墄eM5�֢���
<��+x��ױ�o��|�F��9+*��q�B:��H�N���[?��bXz��G�~��9Xn ��ç�*i6ɳ<�a��X@���g�ګ�����0>:���1�P$�`ȏB!'�16�FCS+:����p
���O��'�k�b��GIB�n愇B!1f���_������]�jh�h��z���\�	�U�gYCx�u��f\�
�Nê��{.ǏU��c�F���߉�[zAhnD���҉��bQ��|buQ7_�\q��0�Y�"
J�`��1���0C�Pt�xÇUomēϯ����QV"(! �0�E�J���N�}�7?u�'�X����>��k��/����4�.�/֑���)3?�SOZ���F4�ƑO!1:�GX�\8�	��/�Z6���L�-����x��klG���<��q�F_s�5���T��[�Y�U�+���S^	<���oQ�|�S:>1�a3�
X��M�#2�I�Ta����cۡ⵪ia5y�%��I����fO%�ⱪ �����*d1\�C*�R(����V��7^����@�`e^�P(��r��e�!ke;�$Z-�&a<W�s���CO��=�(�~�b��EBF�����-�r��>s��'4�_��ׯ���U�ٗ0Q,�pLW�sP�Ž��<����SZp�uĜ�.�F(˒%0�)�2x��ǲQ*�D��?GM]3֬ߌ�����}d��6����� �7, ��Ya�e~I	T�E�# =��f��DC���	\�1
�9�{=�q�:^��������d�Qeԏ3��-LJ,�k�(�J����<i`(�OXJFރ���:�v1��Xq?PH�a�.��������n��(��b�\$�*��3�����d�[��n������Ϯ�P�B��	�x~z,s���˧}�z���y�|�͟�P4u&i�*�r�`������W^���)�z��-0w�HiX
�����k4?�%�����w��_?����S��waR�l/��*��
�2'���H��٫ \B܄5�h�7��j2p� �c�ci��5o,�T�~ǿ@x�J��]��
��܏���Rx�*S_��`�=f5�Vy����{�ڨU�j���碜��o�W_v&�?�`��Y���lz�1`Sۂ՘]��2�Z'I���ڝ��]�c��~h��������H���B�/�����n��z�],�����g�5ʈ-��|�ʗ?��]���f�����|N�(���bQ�,oZW��y��U&wʌx쩧����{���1o��N��i��H��;,r�c%)�E>����E����P���
��e����R����S�Ŏ��JiJF�B�GJfك���EhHn=Ò{`��SJT,�x�1�Se�e�L�%������%���WZ��Z&����A�a��d��}͵�F,B6��/��!���z��4��&E���@>�F$�GѲ��э}G��;������4�6�"��)��_u����מ�n��o���Kol�����^�uh���߀�Ck]@�k�����׾���A!@9a4�#&���,k;�P\Ky�ca��"ʎ����رw/��?�m{�4{	��8�${����#�C��I��RÈ(`	��~�C$d�
�Y*�|Q!+�f�(��9.թp]U��{�`Y�}�G�����(yEh�d]Rՠ�=�^x9��΅��h�_iU�.�O<�4�\&�"���(���
ou�I���� b\�B	!�AD��JԘ=���߀┐�¹5��GJ�2|���`��}�i4�
A�8�$k�4������j���<��md� [�"��VN���)���|��K:Ս�_�����|�G�������~�3�� BJ��\u��H��"�L
!�KbX�`	�y�}�THpJl�%���)ƭ��V�ݏ�y'���ޣ6Xt�ީdq�������x��V����P,�^)�U+X�|R�ق�~�.�pb�&�r�SY���)J���~ =�W�4<���¯�M2M�HX��e��%&�x�|�$�� ��\���gh��r��^	��m�(���$�J7ȽqӘ6�>�����0�=m~���Pl�s &��U��eKe��Z.+ ^���������?��~<��ZgU�4v��A��+N���o|�W'8\V_��mw}����ޑ�\�hQ��a��D]HA[m 7\{�:�d�9(�>���1H��TA�C)	=�݋�|FQNzsKF���{?Ū7��s�r�����~�cګتJ$R9A�Mp�̑�Av��1�|ƅ�g�g�xM�6Q.�aKRS�bh4#ʂ��ҫ���
����{���ǖ�O��¯mc||���*B�y��0�G�Q����P���ɐ��|� 4#�����F���]�0�?��{ueR"�b��BwM���,2�{q�)�_��:���i�4�@H65eG�.,��S������Zq����MAm}������}O��d�@k�L�F~77r�������|���}�g�]��GG�S�%�}pK)��fLn�u�+�/A���EP��)�)�Ix�[.�&
�LO�P*��Q�LM-���ĭ��	��ރ�'�&G�,�R<o�ɐBc�Aq�!��*��(�!�vŅv��|�⠔K�\����bDqM�-���hoCc}����x��������ba����PЄK�-O��	,��n��i [,"�-B��Q�E�Q�30��$��9����8�ezo���0+�;zD1�
�*!q�b��<��@1 `r�dՇ]${wc��F���߃��A��d�����;hhmw�"��:�����CcK;��㻿�~�98�8�'uVS���KO�z��?�'4����ޫ�|��_εz��!�ⳳ�j���k���'�C9��U*�@�A���E�9�K�#
 <WK��8#_41u�t��u'��?Ů���]�hMLnޡA�h�؉���ra�6�Vv���A�M�2I��9������&����;'���	������ש����^镐B�����%#���}���齚��ߏ\6�T*�|��w�b�T�Lers�ꛛa�BH��H�3��Ǿ}ؾ�鼍"9;R7�
�p���vŻ��No��?���D�TDH)#pP;�ڠ�_��{��\+���r�(��J�-�l��K�ĸw4;6(�P�����~�xn�D����C$�a��.^>��o��gNhX���ѕ>���e;iX��H���RF>ُ�(.>�4|�򕰋�
Y�KC��;�+�T����,b3�(����D�9�>�����P�7�}�\�"a�R���%�z�`��C�z���Q�z�BF��OU1����M��fLnk¤��#Aف�V�P 5ш�l�]o��N��H�K�Ī��uTccc��:������1��jlh@m]��ca���C�cO&1<:���ಆ�F466�,%�W�u���s��G"���`�P5�}���1�䢋���4�%�2��
�� �#G�?��y|���n��$Kc��>�U�̫	�Fg`�,m�����ϭz��ѯph �Ǝ���~)��l��E7}����??y�_�x���ù���rWj&r�����ܩ��§nF�pP̥e��l�d�=骧��HC�PS(��>4���X����}�y�OY����P	���� �M��BX�E١A�.�V�,�,�`���"��h��y�j_	!4P�H(oii�k���p�������8z�(҉$��	������9�#k�A�Ecfq�y\F���$�a��niiAW�tvv"^_'��	�3�H�H�QU��F�q����[xs�.�����%�Eja�Vl�`�A��H5�/�4���з'N?i>���/��6�DrT<��.)����C����T(,d�K�,#����E׏�v7�}�Xz���!�DCp�c��L��_��'4�;�}�?=���GF
�X2O��%�v~7���|��k�h�t���k[D͢�8E��"8e|,�pMu��ذe+~�_?���14v/B��e*�6t# ����u��l;)�V��ʧ�+�>m
������������Pu�0��Q��	ط��}�bL��޲Be���BJ[�@�?@,��+�xXCFȫ�@�Ϟ��L8Hfs�
�9��t�XT�-���{*�_��sf���M��\߲���w��h"�Ǝ)h�:�/���`��mxcݻҰ��w�Y��z���j"c�)���ac|�0
�A|��u�
��8�GG
�
�&#E�{�����`��L�D,Z���<����W+2���(:�u5��G`���+�ϸ���O��z䜇�^u���´���R}(���<��"~�8	7\{B~��Q�e[
�$ߊ�.��ᄋGr�^�F��ځ��{���ށU��D����i2�������@%��X��9(v������9�8�E��݉��������ȥRxs��X���=�|6'��H�j
G$;%�V��J7+=D����傌K4�+);�A�N�*B"һ2�0�"����Oc���E�TFM]�Z���=�����ٳ0{�lO�fH��c���K��j�Z�1u�Re���M���&��P��-�(�.��(�{�J�-5��ֆ�|
��v���7�����\�bdx@ԥ+7BM,���]�\���@[{9}��z=~w�ز�6��crd t�� ��X���]7~�������s~��?�ul��6���f~P�U���׾�r	K��!$�F�T�̊;VB�dWT�����D�8�7��z�)M    IDATO=�9^L�>E5�l�㾂��gLVY��>�F65�X؇S����@פ�}
j�!��c��%�ض[6m����0��'�&�PNJ���V)�+�(�EC�s�br6��FF��h�h����ڷ�*�'F�� J�G�c3IR6MH�� �"���$i����2
�2�%S�z���z\p�yX�p>�Ϛ!s`f�8�s����x
-]�:g!r��_߀���OonC6o�uH�`��S���P�[����"�����W���+ܖ|7�? kF
�����de<��s���E�h	E5
%�
�I���!�x�;Փ�x٬���>ub�u�Cg?�ԫw�v3�Z�gXL�)S-�ƊȍbRs=.]yNZ2s�u�T�`l,�\��Kh�\(h��(�ݶ��!�ۼz �x]3l-G�TN&�@,@���.g�M�6�����'cƔ��Ut�� ��-[�z�j�_��R�q�#�`��f�2K(�q��S�{me䯤�Sj��0�LV�%�B��A���xS���ʰ�)y��E�<E�O�/����1#�KJ�`PBr2�A�hʂ._�g��sfτ�q�1<<���b`4���)�9o	�[v��O��]���D��Z����x���(g��ȍ�S��k��I� �>��H�J�`�ĥ����6<���x���� T���V�%Ő��0�T�%�7~��İn��ɳ|�;���O+)8jK ����%(Na�A&9�,�Yq�<,_�-�m�ʖ-�T�B����~��n��>:_$�`$E�� �/	����b#�A},�%�f`���X�`�0sj'� �z�5<���8���lz#��|����,��}K-M�,4�j�x����w
��<�ٌP��y�Oz �p� �b4��a���T2�\.�������35╆���O�?'��PP0-�M�b	V��p0��sf�ܳ��ҥKaĢ�{z��i�v�&Ә6{�Ϟ�t���|o�s{���B��4G�f>�SBzl ��Cįa�N�yƩ��Q�F����a��Cر}7�������Mp|5�+~��8��_+#���/��;_���Y�~��{z����� q�D�墸X�z��'FG`(��q��ڌ��.��O�I&�k�m>|�w����(J�b�t�X-E�="E�AX8w*ϛ�y3���T���m�]�e�z<��c8�?B�0Q�u��qL�������4uXV�!�`?�q4�`m�;ﴷ���l�F9I�/��wT�Լp*������nttC��$�e�q�(�H��b��x��}���jj0�Hc<�A>_��@�P,�fL��SO�i+V��c��hG��֭�%�]�x1:��������Ko`ûېΖ�+�0ˎtIX9a�q>	+��$��	c�\D,�,���6ؗ���A��ʖ�Z�]y*U�<���!PܠFR-������G=a(���ז�����z{����Ѱ��/�>�K�^a�f�H'F��9(�)x� ��pB`��Y+���jz�f�>�Pl��0�tMnǩ��ӖaRS-�~p?�{s5�X��ݏ�HT<��mI�W|v��1%���˶t��A�DwO�����'O�ܹs1g�\455�����N�ou��f4&���jÄ�U=�D�#X��^o^��)�<�E6�e��Ç��{��8�\�BV�����92:�d&�u3:r�4�,^��\r��uK���tdd��Y�P�KN;�x����S/�®��Hd��ґ����P���.�-�G�$�Ơ���&�/"�A,������Ï���L��B�v`Y���.����.X�}�w����OhX�>�������o�8��T�p���^)�b#���S�cq�V�����k�^��M�	�$�p�s��bq١��`@C,P��p�%+1��N���_����x�'p��>4���'����̬��G��ދ,=��D&#�r��N}��gbj�4�[0_~���1��+u�b!_�v^����I�����G0S%L�А�KC�����
&��=^�l	���\s9���b߾}
��L	����H��/� );��Y�T��9�p�ޏ�3<�9�7֬��1u*&O[��T	y�y��z
�������$ۖV1�=F�Jy�:RXP��1J��c���2�(��TTX�r�8�V*}�)�o��?��?�X����cw����"G��т���R�'�e��{�����}���L*��E~�A��p($��X �(B��BLJy�M��^}��8��˅<ʙ�nڌ�o�E<��-�q�P�F��>OJ��R&��qCa�uv`�i+�줓oh���#�ϡP6���#G㢄�!�.p�����b��.�|b��R���碁�s����~?,fX���� �-�"����4߱3HlܹG����1�&�)�<�����iT��oļq��+��܌P؏;�Ɔ���6O:NЏ����_~
�C	i�Q}>�39)��P9�l� !V�2��F�pe8��_�Y�fњR�$�%��Q/�eV�2�����zb��؋��y������[D�e+j1)Kc�k�Z��j+�t���z�.��X<f}P%d�5��c���5,]:�\t��.� W?�ك�|Zxڔ.u�A~+/�1�ҹb�h�hLąL��� �M����?_HH-Fzt��Ò�W�8. �`U:\[[#��j?��=5�Va�ӞT�gMT6N����76��L��j8�7%=�����E���b��s�Q`b��H������+���>44 �&J���
��\�ꐋ.�_z1Ԁ��!�ر}��X�l�gvb�$���3X�qJ��<;�?�E��q�)
��"�5��Q�
�"���rv�1� 	!�L�g/:��S?��-��S���#�ܹmw�������c��ɵ�������rOo��X[I�E�P�j���)���X�RӦ4a񂙸��s�O�"=6�Lb{v����0Z����^|����K��
崛��QY���V�u��8��h�4	f���G��Ho��|z
��4(d!M�>�B__�`���8p@�����蛙�z���L6-���4Nx4��o�y��`����>�[�_MM�x�j�H�4X�e�D�X�r�X���E��hZ��e\���Ƒ#�P���`hD���)x��5`�Ÿ���Q�P�T2��w��o �͓�`�)�4௏����=��TIdŅ=`P >�7��i��.E���9ej�t]朸Y�>T<�g##�L�e/X:��?����=�a�����~��;v�8�K*bH�j���׺Ms~G����D�A��)B��@wY�rq��sq��Kp����4��9�l��&�U��4��0DC!�c��H<Z;&��s����K������ ��چz��5^�&���ڵkqp�Y8�z���3<P�P߄p�e�	��\F��H�䤳��vtt］���&�!�،s@o8c�̟?_�輹s+�!�z4j�T5���3y��I�BO���O`hx c�	���4���^�8����م}�z�[8_��{����͛��`��%��5��u�H�]�P�Z���2UhR�e�4����0D^�
���oH�ұ��W�h�H�T���'_�ğOhX~��y�������?�oK
����h�l����D;e��3i���Gf|P'?���PFߑCȥ���s�c"P9�Ch�R�X�+	K��
hlj�y+/���]*�o����GG�3M�-���0�c8t�V�Z�6�����p��.��g����*��u�\�$�^.S?���;Y�v�3�j�,.^S'!%96.�κ"���Ja����k��JBap\]]]�5k�d��cⵘ�UN	d���ey_c[���R&#�߶m��~�fc�q���
f2Ԁx�K��篼Z@G�`/֭_WW�O���ï~{I!mG*�J6T�Y.հ<��;��h���kIq��DԨyYdհ�����:>��_���'�XO�:����;{�(�A	���a_y�����*�����Į^=�Y�D?fO��_�>�Dسu+�:�H �|2�0�������S*��#bd|�P@ ��W^��I8|�0>$�P˅o P�ū���Kxꩧ�}�N�C~�~����+q�I'Ix��!.�岰��!h��XW�w�Qѫ44�y*��LYv��,0 �g*��tm{�@z���u���o͚5ؽ{�������'�,*�Ky��<Fo������B��y��޽{��ؽs7���(�Eq�'?�9��A���o\�C�c�%X��4���0����8p8%��i��f���VIN@��4V|>Xf�cUd5��`�=��d��:?�/}��'4��}y���=�����=���Q1,����~��N)���ܖM�y��[F9;��������-AH���O!3>�cAD����fYR�#Hw5ea�Kh�.��.A&����;���YLN<�A��C�����Z%��sΑ��`�"YH�%�ᄋ���Ѱ_~|<)a��Df\k��P����Zb����4B���dѝ��k�M�@td���?ϰƐ��~$c�)�=�\9��^����Li��m���"$gs���/�4�A� ���������}�^�H$�t&��7`pp��]8�q���_���x{�Q�]?�G7P�J��Zl\����o�d�J���0VM8�H8�r�������+��?5���y�����;����y,�	�E�X�\�E<�'��\XVٙ!�<,$?��fcJk->r�e���xk�K(d��BR�SY�������@�
�4⍍8��Xq��D�8t�06n~[�xS:��y�B��f5{�1�WK�-Ź�'$hcK�`+�h<]�h��^�����Oג0�	����FU�"�ez@5A�\��Z ;�=0OH�Vտ�fU@�p�5y𻪽���K�W�¶��J�@]��,Y�X<^!�fᒈݚPW_/�:�S����b�w@�h���Y眉�߷-�R;$�w�!�N�Ɗ����#)��Ď�H�A���T��Q�ʶ�wO�S���3�j�X(�p(�r�Ͼxy����>���/Ϲ��'o{{W�y���y���ҰH9T���aI{���ǲ�R�#������/�"��>��Ckst��8uO.��[Md7d����KK����*e���}���j�{�4���ׯ���ߏ#�	P��5������O�Ԡ^&�E���������%؜I6�{r���xD�d�YL횂t6%\��,'�
y���H8�\X������r��$i���q$��f�BW0�Ҡ��[�7nƮ�{0�{�:�l45���Lf���(����"��ql��c�ƍ�Je�ܽ���*(j/��b4��
��a��?tS���¥Kq���y�y��q7�.�+\9K���k@�xK`�jK�E�1
��Q�u/\��՟��ɟ�а~�Y�>���_߸g��G���E8�_Կ�
9�a|~]p��`("hMȇ|jN)�����K/@>9��xM��&(&uL���D,��~�%���514��K�Grs��w�n�&Y��
��a�z�{�ط� .��b���Wc��i2�@#c�ӣ�1 .��5M��Y��Q.B�S���>4��c��
V��#��9IԔ�"�l�*���Eb4!)Ho]9�N�fIj�^g����^J���ՌP�*�hJ�Y�ڸn��X��%D2�d�"�뎧hkoA[[;̊���5���~�� ݐO"�)���I���;m߽�6mY3�b�
�'���=���U���a9&�#��5G���$S�1
0x���HAM(���!�������g����Wg>�ȋ?]�q�����F%�0�sHmS$)�dة��Osa����c��)����3x��Q#���"H,�V�k��aԠ��~,;�T)��a,���w�"A��/�];w���\}��v"_*���=�����_�I�-�P�G�;�����Wh������G:�����C �k��1�W�D
��=�X8$����H7��=�kʔ)"?�7�6���+h�4.�Ħ�	��$۴�heaŏ���zbٲe⑉e��ƒ�2~6�̙3GX|��߽���B	C�O�102�����O|\�b����oaϮmX0�-;{�˸��'�«k�h5P}up�����(I��cD7Oâ׎j�:��'�����NhX�>���{{��ol�{�W�����M�Ov��2�VNlg�e#�3�(�I`��N\��K�\��u� "��d��LN��f\lL�����uL�"*�d6���Q����c�d�n��v�>���b��R�܅�����Z'.P(��#�	�Zhhcc#"�,\4��앾��I��־�^`ɒe��k׾!�������`/�7z�����Q�u1,�3���Z��@�0����G���1��T5Tx�$K^Oc8*�(�K�i��x����{� ���j	��#C��H�P�2}�l|~2i9**�t*�����A����p:�LA}S�W�~���A��y�u�Yxw� �{�Yl|{/2%%ǀ���T��o���(�"��H��E�'}�o�{'6��_�q����M{�,�/�z,!;���!��12������.@1=���q�uW�ʎ��'�����
�l�e���Y�s�?\r$��<O"sn���a��i⁞y�Y���K�:u*>�яb�ȥ�	�#�6+�
K$1}�t��w@���v�V�£�>��o�Y����3�bQ,�;O8���1��O;]0�`� f͙-�;�E>�EK[3jk����C(yqb,���Ai�hnn����o7��Cԡ�g��c9����|B��h�t�+�T:fh��P����9�D���;o�,_&~z=�A�`(&!
������X��-�,��z���/�r����_/��r�uo�!�7s�)X�t1^]�w��f1��Q�O2Q��/}�%p�ʍ0=V0���~\���[�}��'6��^\7�O>~��-�W��/$M�rԳS�}�+]��t
55qhv	��^i=���>�-�G�*:�����X(,��J�K�+�t�gCCC��s>ؽ�İ�䓑H&�K�ܵ�f��g?�Y��FF��OL�Ѐ�1�����n�֭����*�s�n��3gΔש8hni��f �C*��F/3"Jr2���/y"�}����(�:ڤ�י���u"ʣGd��?�z�@�͛'��;�#t��%X��$�	���"�180,?s��rU�3���
��Q9�hАv�ޅI����+���%).3,O`�E�^z	���yO&�w�A�L+W�ĥ�\&<�-`Ӗ�ؼu.���hh������<���,�Y�/�	xg����%x��K۾��o}�'�Xϼ�~Ɲ�?��uo� �CA�a9���%<�]�d��5��1Ĵ,>����&ּ�J�q4Մ���)r��9W<q��6�Ț:��x}���锰�S�����6o�/� ���O?�\r��7b%���&lv}��h8+W�O�m�wkk�t�݋��{�*��SO>IvߪW_/Hp�H��Ȝ�=S&wJ����N�lG[K3�z���Z�f�M'SR����*��14r�ɐO�:E2�ށA���P����ċ�VY�'���"��V����]�њ���4�H��[>)�mxlTB%=3=WM��b��|[6oDmmT67��� >r�G�x�"qܷ[�y��c����#�Ҁ;�{���C��Xz�/&ԓ�6?��I�4�CM,���!�3����/~�����kkg����~���C�MUt���Q�bA�}��lVn:�ɢ�������g����y��z3�&�%�S�� �rA�m���/ �XM|����R��J\���ױn��u�9������$�L���k||S�uc۶�R�8���er��G�d������kV��?w�x�Tr�W�Cڲe�����F�V9tX��J-o1�\!'!�m\�i8x� A@��mm�G��    IDAT"��S�JH������-����ӲI��ldxL*�lU� �7q,�E����{��!����x;��믿�j�!��l�𡵕�����lz;����38��t��`΂%pM=�I٫a�$�~�E�3f����zz5�-3`�[�a���	%m�ш��?��qμ���_��	��՛g�q�ÿݰ��Yi4$�����&�|:�xM*O.�!ݼi���g?��k^³O>���Lii��
��O�,�4z?�ı?�tu4�t�t�`���%���ػw.��2�{�����,�A��Ԟ=���6i�$������ŋq�Yg�'��]?g���54(rWlL%�Z��b�&��� ���q����F�%�m���X]�����b��`�CK����#�#OE�ZU7�癳���ٳWd���f`��S�m�v��� 0Q�=RE���k0T�p��64
�B0�!��6����w���`%����FM���M��;n�`�Q46�K��h���?t���5orc���u������o<����s�E;a�q�h+�TJ���gOt�G��9���������Ϯ�󗇞���v�aRV��T:fI
&��+�TR#0�<���_An�0���m�	�1c�T�����u�S_(gU}�0�<���E���u#�$f̙!���^���.�y�'���^��4M�04����+���mܴ	���5�;�m���1�[�3�֦f,X8O01
�sb3.>K*���!���/Ac�g�"�`�dur�\�m���ر�{˦hii����I�m�I�<c�l>e<�����0m�L�ٻ�<���I���X�Ḉ���x���:ሧ�%>�����}�qL�~��O"����˦tM����?��;��KᝆJ�\�`��ȇkl�o���^}�%|�ӟFیY��o���Q���Ht9S�2������J�bYw��������֓�o�{�}O���-{VXi>Z��ݢ�:�j>�Bvl v)�/�&t���Ϸ߆|rs�MG]$�Ȟ@:���&A�܂�d��φQ�w��hnm�c�xk�:q��\s�����p8�\hb$���
�NP{�i���܋��f\x�y�N ��i�,��~��5�EN���9�\��˗�B���HV��b25.N�/
R�@o��@�بX��Hw�-���(r��)
T���O�8��<f��1<|�G�g�y*ּ�vn�*uɖ�6�Hof���� �0:<(��^K�U�3���=^Q���n�,�㤁rNn�çc˦�x��'�ͤ�t�"�	���)g���/��Dr �U/��ޞ�����#>���������QP�P3��V	-�qDI���i��~r�O��o'�X/��s����w���u��A�������;���Ǌes��ƋO?�7_}3�:���$�[2�Պ���~�eR�c���QJ�'wtJid�ַ�?��+��N�e
.6a8� �K�'	�������6lX���8�#�"�e��[k�b||3���.?|���뮻N�,�4"z��_;w�D�6&��顣��_�X�v�B&�Ŕ)]�1�D���"���kr��4���4\���'��O�O��k�41����ªW�ż��q�+1::.z+~�FJ:�ܘ���#�A�tNő#=bd�-��� ~�Qy����%�ir�E|� �twU�v����ȦS%h����ӟĴ�s�����.֭}��;q�Eb�����߇�G�pH缺p}MDHqd�tj��w��_>�a��ڦY����;ֽ�o����fBv6���s9��D4���g1ڷ��ט�T���6)B�� �4�퍥R�<a���R6���t��{�ʋ��,E�J#����W�Vlܸ��8/����K����?'����O�#0]�t��j�06m\�1�Sp�h�xA��1�������V�^�:�K���.�۩�

@f�u`��jąR\��OΜ����u-�hƒPmm-26��L>�DrsfN���������8���+IHF�}׮����<wA�e�z{�Ż644	I������^��r�`7n4z��I�P�� �P��o�-v�؉��z1����
h���0�k&�cI���j<ڃ�.��3�q۟��_�|��Wg��!���懱������׭_8�a����_���?Ѱ,��;[�����h��"9������K�M��o�1P�cJ[#�"a�%vL�K74���p��E�����$ڼ�m���/©+N���ޙt��XS���pR���%�����Уq���@��W�p]t�,doO�Ϝ�ɓ���عS&�!&���-��ၜӶm;� �'mo�@���4"f��X�V��Y����܈�Gze̓�P!����NMMLj��tRZ��餌� }ƌn�l߾ﾻg�q6.��J�zm�����8�Ν#�7��^���z-O[;�E���?���}۷o�@�6�e ���CR�eҒؐ>ٸ�\z��Xy��(�8|�(�X���c�Wc(U¯��w��1bHel�19B2ѿ�'�~�ǟ}�s'4���ޞ��_�uφ��[��u�OJ
��J�,�щ�}�Sx����W1�����-��.���5����L&�
!������[ZZ�¥P
--�^h���P�X	�ɸ����3���%<������9s����^���R��B�K�ƼՋK�Ago<}�D�% ��b�Ħ-�����H#���,��=o!sVw<̣��������)��a�"��B<���F����ILL�('��cb%3Dt}rf�!�J�)rRQQ�̌Uz-�DD�}���/{/\���h.U�d�rh����<���nkk�����/>^�����J����s�D>JJ���ko���F1�}�,�	�����Y�2Q�ufv^��Q12�^x��s�΄����I!��g�䄊�B���K�����7j��oAxx$FF'Q]ׄ��Zħ�!u�*TԷ�7?AAE+-]a��	wL�t"�������yY����<�ɧ����#k��I+�ԡ_Y����1���Af\���o�
Sc�n� �H�����YZYa�lFsG�]�%�J�����d�(�6`M�j������F64h҃�����#F�D�u��1StD��P�x&�}�J��hh�q�F>6���*DG� 3+KU]W+��|�R���Ɣ��$��Dn#K������z}�_��U����ފ��j����s���Fn���.hjjVe�����Ҵ�����)X(p���N�hB�aQ��mĐiTy��k�C}}-����	��J���٦P�pNw�wU��v}V�%%%��w�����ަ3$Յ��Q��^{��92����wKIO��������;zP^Y���N�߲i���������¼���\��o97�$���_���z��<�����9��h��շ˳��CNb$���o����CZb"���<;�)�n
�*&���2j���֬�l�
�qL�o��f8�;cz�ފ�cF˃9
���1�S�u<Ē�by5V:
K+��%�A� '4��U�V���O�l�����O�4Jug��{��&��jj���o��F$�H�j~nA�͖
{�mc����H�����Qsc-��twSh�B����S��������`��<�024 7Wx{Rsu	�~��56�`rr�v����O>�XƐ�*gϟQ#��ތ����n�l�g�ux��uIk���eX4>&�|���_��Ձ��,�B�]��[�����bϜ;��y3n��0�Z�7xu퓘�r�� F�Z��g���~��u�Le��x�����us����ъV;
�������<��#64H`��"��k��"��-�%�Cɠ�I3||�������_��H E����u�q�YaW�V�G#a�����X�f��B�������cH���S����ũ���ގ�^+��Z���R��s�x��ShXʵ�����^��8���&9�ބ7>6.Z�sUe9RҒ���Pq�x��!-)E�Alx����z�ċ�����B8��r����N��%�P�ڣ�1	� �G^Vu]�.�m�݆s�O�7^ŭ�ތ�o�V�����չ�������N��|��q���۷O�/1�=���3J���쟞� �*
��u~W\y���Ҋ��&���c��ݰ��{�.���]E�w���>���
OUD���7^.�n�0�l-z*�8�ؾ.߻� ^���h�*GBd8}}/PnG@�?`����ƶv�xxb�<_?���*̕�2`�>d2I�wf��{���a����ĲX�������a1��5�����nkc��ή.���8qB�h'W_+��/����\�?�#2#�'Ҏ����� �^�dT�frj֖�v�02jR���\~��d��IMMEdL��2%�2�!�VWS��0+3�M����
�������F`yy�>��vx}����\wõ�����(<r�&'�e͐Nb:�|�Tί��
���?��;��xv�.P�����Gﾋ5�W���#�j��HM�F[Kf��q��rw�Ǐ1<��P�>�9g̎ �g�/����'����?�x���i��²��u,O�ే���WhO��D !*B�$}qښ9]�� GF��Iqeh!�Hj/E�֯_����-̋��ǜ���U�����~BW�����`_�Ƭ�������g�oº��e$
_~�U\����ގ!6П��@,_cjr�^^�:��1L[�f�+JE�KL�CNN��pxdP-!�&fV�ͽ��1��k�76��t����}�#W���ũ����vRZ*��Q��7W/�|2^	O6�e<w�rsW#7wN�<�j������c��m��a�4����s1X�̳�ax���Q*B"��W��3�-:��C]S3�lށ�W_���4Їޞvy�m�����W���+���S�_���$����y�����ȉ����7������t����k3����܂���VW!+%~^������PvN�8y��t�풅�Y\����ض�V1���jy22y��8��0H$����"8肊���'�y�M�33hhh����1���2���D?V�4l~�E4l2��w�o���c�����d�֤_���n���nh��6�#�<������C��GV�*M�����#2/b8b!@��7'�Y4�ՋV̋�;Ї��Aц8���V�LΙ�U�T��ɟw��q]V����"���)&~����%�*�BB(w�q����7���I'����Ly��>��>�k�����޽����2ѮY�L�q�~��W���/��u�����3�<���։�O���7�j[��-s$k3�x�gw�ay����	�+��R0�ע�����Z��74
w_��(�L������+U�[V`�6�f�"=nV���ب$��*4,6���R���|(z���H����Ao�PnX���h�m�`�**���h�ԩ���r1�fx�322r�'�cغu���а	��~�Y��ަ�457���Q�i��uP����SF�<��?_����_�G����W�m�U~�)�4�5kV��O�"11N�;?3�cY�������x�8~����y�����g���r��Y����������^�xx���^��<�����ۃ�C��Ԟ�{����/>h2��3�}�Z�dd�o�±�����@T����>��m� ����W��-�|�W_.���>����A�9�����g/`uZ<�	�17gVn��ggW���� �2BLd�-E�ɞ����:cc#�V�62,z�I���Ј�t&��-�2C;~CÃ�H|-z���~����T=������N-S^A�6�������kd|U�uW�(�bϒ�M��V<X�"ٴy#:�;p��Y�τ�4�X;���S\�-[6)�^8����� UUpuq��#�gϞGum֮˃��;L������Ȳ����**�%�rTVT�7bDeؽ{�Ό�)��(���{��wߍ��6*�����epdHn �y�����܉1==���r�	�DIA�]>;�9��\p��Gk����{�)"��z�Ƿ|+))���_}mX�˻��~��WN�l�_���� ��z��������6�N�T賴X���0�`c� [;{�uucdrsǶ��!���[�!0�O�Ź�e�%����..Y�
.��^�
�Ř����
C��4�97'�����Mh�,�)���7�Th۱c�0*�J�B��ID�D���5u�YZ���7��k��mbcc��ҳ1�fu��RSC��G����ș�$de�[Ц�����$>^^��o���"�c���ҒrQ�SR����Jy6��<<�����s��]����b�w��(�P�/OGFv���:Z�18%C�=Xll���J��3��=��fx�T싋�Ab|�"�ݩ�'��� fĶm۰:o#:Z�0:>���*�����nE|R2^x�$>��|�,����zG|������%�_x�S�ֲ?h������7��.�_�|�S�4ljoe'$����ZۉS���G�FG&*]rnn�l� J	F�3�X�sF�������]d�&���0_1��V��I8 �����N�|}�''�I���c��U⎕��`uvr�rP\\7QyH�������S6+�4tVi���J��C���X�j��de���$��8���Mbk11hok��a/O�GF���
�����h�������Gl��iŦ�y��4�t544ay�R�olL�t��"BQ�X���y[N��S��F��D޺�����%l���R���'23ӵۨ�\>^~��XX��� ��s�������d��s���5�^��
���Sp���������	���hX�eu�O����O�:��׹iɸ��o����=����HW~�47'[{i	8��`��u--R�[���a�\�+f�+=#U��yl\	&>���� U6h����5L@#���S3u͚��d7���NU@p�@��.�;`���
��~��+:*}�T���]����C�<o%�oek�U��1=����N�Olذnn.ʟ�ڄ�;66���M�0q�qwv��ܹ3��O��*G��^쭵��X@�@�B�yb[,���B������4+OsŇF��ٮA���Hc�X�ӬF?��cl޴�ٹx��wa�U�;�H�g�nTT�!5%I�pa	�W=�}�գ��c���r9�b�K�̔�}�'��Xaإ�
AYY�(P�7XX���f
>෿{���C����;��↾ѰNU�G<�����Ͽ�j��?��[HO��o~q�և�ƅ�#�aGk[XP@��C�sh�hWÖ��ia�6� ^�����ޮ����e�Ɵ9#���a>�6�aa���QC"�<���[��2��0?�<�:����$FDcc���+V�HNID�_8Ξ��z�������V���eJN׮�ASs3j�09ŉhkxz�����U(nV]U��tLL�B���r�6YT8�yK|���i�)�qS]M �.�NF��Cؙ���4"��3\1�rw���بZST.��--.���J�Pjz���#c�r��FeE� ��n�1Qb�::p��cv��%�f^�������)�UV��Hb���h�px��q���r2�شe�<)/F���:;��DVN:�|�=�~t׷o�vjj��7VAE}����;���禦���CѩSx��W����,9X�c�d�205���n}@2�<��T�tJZz���p�cE���!zƸ�f5�nۺ�<������L����088HK�<{X�a!AXE��13M�ppr��=[P�P�sg�0=5��B����`||ˋ����CdTZ[)�1����خ���M���R��z(��t�3�yH[���L�(mD�d��6w�&��u��3�f����|44�)�f�oCYY�*�uyk%��"���[xSss�*Wj�3g=~�$~xFW�    IDAT�=ʛ��y�s��b׮���<aool��a�H��W.���>'\����kQ`:�Ĕ$t����w�Fu��k�*ޱk���Ҳ
�9�����߄��:|���o�ᚻ���s�UX��������Ϗe�$$�����=� �F����yq�YQU�z�RlЖ�~�������&WpŕW�`�i���'̪�X�WF6%�NF����ё!DE�&�ޯʆM�Ӡ����v�ns3ӘGsS�&�3W�����.`jr7\��|���?{Y9�����r��u!<"X!L���l9|���j���}�����΂bhhPF�m�feYy����s ����D�3�����N��L��Ќ�{\��N�/<,D!����Ξ���<|��$�K��_`�J~�b���| �Q�K�[|��n�e��2� nF�ܡ��'��⩐��?^R������\����>����Ȉ�1fd�p�\�����Ÿ����g{��w^�|���C����*�PV�����C�g���;��'~�����r��ҼT��Yl-m`C�eg�ڶN�&�S>���D�P�A�X�a�p)~8��ı��z z2�ff��;:8Ї�W쓞B[sff��P�_���#c#b�rp���)��DYu%�-�����~�D'qg(rqv�7ތʊ:t��b�b7�x�ͣ(/)������^�������#g��ϧ�z�_=��]��U�Sb�(Ǻ�fU�q_-Vg���N�=1�А@tv�ctlX�0@]]�[��慭[v���M�x�GƐ�6���X%����@��8rTޛ��vK/ગ��EY%�X���*���oN�jU����Rh�,�|�|��ւ�����L<���F�<�i2/�ةSg�c�n�o����9�i?�l(,���}��?�q����'�-JΟ�o�����p�
[+n�\������x�cS�h3a�,��%D�DX�&W�� �9ˊ�骷W�E�&'j2�����P��J]eƌ��0!�t���2Μ�\��Gp�w �v�P�`m+�#�&8���VYu��������WN�>�ə��~FeY!�|<U0�L�
E�Ѻ#�F�H�>"2�+��V�'� =#�C}R�����������_`&1'�'^oo��9arju5���ԐnAA�<��_""cT����#:.V���"A@�/*�K�������|��ԧ����ٴ7$%-!��%��O>�۶�s���IxeݦX��ŋ/��Ç�ܯ��2<xc_�)�I�ﳣ_ 6!��֭�N�y�����yyy#�豪���~q��ouuu�<��/�'���Z��ɒ<Qv��k[���6�����{lL�p�.�=Û�s�n��K4s+Q���_bQ,�	����_��\_O��f�g�V�pH���<<<�q@�b���:��� 45����K4;[%�darB��Rw����;gAaek����,� '+S-�O?=���-X�nŃ����x���ccCjwq��^���S%o���8�=00���lUT�q�UvV||<QW[���͛6���Z�+<2�1q� ��7 /���>�^��Q4��|<=ĳ��!Nu錸����K�;1>~��M�E��O»ﾋ��=K���lAm۾U
������Ι��mߺC��pjfU�5:��|�Ns�@�O'�������fê��z�G߲��ȹ妛��}?���%�c�a����Yႇ�I^n> �>JM���J?_%�4*Vz�
���vZ���vL��o�C�bQeJ�twu��؎��HJJ@O�1X@Dzժ�zH�-��6'��ͮ}Ww�򺤔dx��(w��g#���G?="Ȃe�<� �t2zU�M��Iu���l(��P���.񵄄x{UUr�0�9��< Ʌ���� #1���P�$�G؅�Vsc�����p#V���Zm� ��ʺ��Tjun.F�F4�A�%z$
�0���tv��ǰ:7O�Ӡ�_���O�����x)B�,�,�yQ���P��gGT�S��C'�n�
��E�e8$i0.!Y�#��M�����t���?&FG�_y���}���Z���G:ȣ��2Ӓ���,����s�6O����1y�q�A�r���(�.�_q��h�t|B� �g�Bf&�����Dz�qS�W�E��/�/���D41!Y���CV�+q:X���9U���M�kh�!#5$( �M���r�k�N��u3��;:9�LLHR��y��Nxyy�3�p@�};�"O/7y*bT�^���H�������_�R}�G�g0)���P���\���Ubp���!1)M�â���!;'����7cvnʘ(��R��OP��9I��8��H��eJ�7��2�8a1��s0=ׅ�jk}��g�2���Y$1�!7��#�?������j�ؗ'T��ݵsgSrR�.{{����[���n�TUU�<��G_ٶm���&����X��7,LO�Z��H?�F�Ʉ��E8�{���������AÑN�ܜ�t�t�����ʪr�n���#��%���|0'O���XhX�$���5�<19���PlشU�U2`np��`eYSY!�۶����#4t�&(Bjoq_ǯ1����6�*����`��"-..DcS�4N��W��y ��	��YX�(�ڢ�҈�w�g��"���+ݫ��RQWXuI����X��
�N�8u��:�����bb|R ���� ��yy�#h�lW�Ix�a���)az���w�C���E8�b�*]��c��y��b�p/6���1��|���?qJ�mjiE\||��7:::v]ְ***��~�/�����_zE�v�*8X��qXrۻ���m����jpb����߈�EP����1�oL�d����v�>���Nxx�*#6}*;��|��D�痱e�vi4���KX�z&g'��R����ڡ�`�916���x�Y��҂"!�Y٩J�	Q�:s�7mEZF&�q��IDG����S��@hcc- �a�?yb6V������bb�����)~ӎ�[������Y�Q���Jy���7J#���H!��T
m��u`��������qM��%(B��8��X,c�0'��c�y)���*tjC���rp��?0H�v�4ll˘�����!�B(��WTP��_~Y�yN����;��|y�l���2R.]��m����]wYê����ٿ�}Ǯ����C�%&���bs��\\�{��%Yh��G���R�040�\��+�4v�P���5~h
���Ò���"����)������k��ZD=����fM��4�;N������݅cǏ`|bN�N�b��0O.���NOᖛ�G{SN;['Q}�2���R�ƆV1��h�<g�h 99�u��81�۲u��l�o0�Z�v�>�]�}������a\�p�\�����L��2.=���x���DANz���P�ڽ55�������-�Ӓ`�@ͭ^C�"!�E�������������/u$���?b��+�n`��Ϥg��]n�$�����0��j�މ����s�������><��38��g����(�>q�
)N�[ZZ��رc����۰<����c"co{������ђkp�a��"�-�uga���.�&F�OЅ�(����xx�i`�v�t��Ri�P��y��W�c�,����m����,��	���܀�ɑ�ʊb�����U�s��(����4�7!%)M�aGW�0�͛��' ���]�j04j|�P9H��MMM�1�W��uk�"8$�!z�-͍
���45��j�PN����'��¾}���ت�B��+�3g�ا���rD�#UiXA!�8�[�R�[��;"ʐ����؈�{��e�#�3/"�[|�$D�@X�ѰB�#��;�H�I;�,�Uʯ��/�+������_�R�dEE���kfffd�����GGn� Ҋ�
���҇&���=����==\a�e�s󰳴�ȄG�؛���D8�[�v��E,������bb�
�����᭢c������3Vc�3.��u~�/��,WM��;+�,�oh1��B��;��b�
���w���8�8b�ޫPPR&��޽���~9yM�
Ë��=��Tb|l
k�6H����M�>.;�
�I�J{�ǑT�ih�l쇒���ֶN��#)!�܋��B�T�"48��	2��V�z�M�Z����#vn�W<٫r�/�U�����Da����_ɒ���~%Ʉ����������OL7����ܬ,�]�r�w�|/���"��~�3!�M*��������طg�S�b�__'�'N���5��8�ũg_{�۴�T��ZaynZ[����5jei�љY4��ch|!��:���£a\���2�,쿆h�L��&��6�U"C��փ�{�67��T�М���s�v45�kގyBvV:F�{P\t�n\�{XX�cj�|�����w �b����������Ҳj�"{�*��y(����׍%��GLę���0K[LO�#(0�	ih�hFUm	�]l���%����W���iz��X��
Y=�Z�	;KL�����
!A�HMJ�`� Ξ����(U��!(()���7���11=���a\��#&���c�E
ϕgJ��%s+A
�˂d.E^�����T� EhY�������g�v�9���{Ժ�4 ���_QU	�W�������������#Gnx���^���g��k�5�M��%���Z���7:��	�c�HMC_o�n
×�@++�QL��%y+> �"9A,�tZBzO�vl�£��D'���ˋ8�N��LNsWe����:q�9���0W���˨�b�ηp�d����Ľ���}�������!�I�����#g���@��W"P[TX,�@_� 5�	�.,��?�#c}������P���!VN���Rȗ"��jI�E��2���T�����c]�z��V`dpNnؽ�
TU֪��
��������"a���FlZ��q6���i������f_Q�D:{�@/_��'&e�����A@g@�RDd�H��>�,���q�=?���Ey�y���e��s|����wDEE}3@����W��O���P���ٔ��*^+�p(�
]}����|)s����Lf��e��[�7KCo�����[���o���m��~^0�r=G Ɔ��kٙYHN�GA�y1W�=��X��ioQ���%�8���73;�^����^w#�����
++��݀����6�"�HK�"tsc�g&01>�x�+���k��c��r���Լ�P!!~HM���� jj���Pgx/*(AhH���}�C8s����i�S3�(�(���=��\aog�ٙE���?�b���WU����)iZ�YXV$(cǮ�}s�aBl��ҝ=}�kegr�(_����D�T��6�*��k�P��0��/<��5�\c, ���gt�n��v�ڻG��9с�f����mc��X}����?��+Ã�α�Ѱ��Ԋr�����-.[����Ұ"���١P�C����Qj��=? C�[;�vİ�`[i���a��=�7�������?x�gf�Zm��l����������#�cb�9p��Y�Lϋ�@����a��?g訏����5��F|\*6m�%o��ӊ�zU�ӓf�<��}ܱo�^u��K�jd�ujH�`av��~��Z��H&��5�HO�u$}�2�#>!I��h�oS�F��hko������uy�-M�Q�nڸ�����F������휜���韛hݝ]J��6����9�]X����dm�%k�g�aX6^�~5��?���|�%�Er L�9Q�v�F���Ȱx񹈀ޜv�駟J6������/���ƛӢ�������߿��;~���^�Ĳs��P�dr�6��kv~Y2�����S�Ƕ
=8~ �j�d�	�F"��B��&���1�d���~���=��ۄ:heL/�P���*�$�j��\-��n������3�fRv[�[V���|������td���yb�U2a��՘��4�e#��Ī��˕�{Pp(J��099��k7"""
U���EZj�0*��L�`��XY�FQq%f�V$$����X-���Y-2���#zJWg����ظx%Ԥ s��$�h8/@f*ϔ�s3�X�R�Ғ/�T�Ֆ����E��w�vR��Mt���𧇌�Ass��o߱CFM��=W\)��s����Zj��56��֝߾muZZ�e�7�8��x������e�%щ�O�I�u�g��Ձ	���D���Ӈ�n�d���5�����d�����ݻw����g4�05e�C���M���N+=��SJ��C�EF�<5/(='�q>���RlڼA�S3<�{w/�[�	�N�Q-.:nھ�j�LʈP����Ԃ����Ǉ�[)��n�:Cnk��̴�#��H�IH���1-W�����0� 3+Ed<�҆���������2��2�`�C˓���F�l+� $,X^Z.e�{��p����b;q⸚�T�fo�?�H?��P�Isr�hX4��'��y����\�́��{�1�l�!��Es2��&��|A�;n�����W7^ְ^���z����]�ÂB��8'��	)�q[����S�pvw����Ձ�`�;шHd�~i;֥Ig�bX�����7v����#F<�ȧ�F�x��AyI-����c�@%�<z��+�S�l��wv
͍����j*��qEN��ٳ��'%$�������9��$�%����#)%M8�[����$�^����⬬x�ڣ��	����M;1a������@BR"�Z����K��WI��b�)I/����`��5��^��|K����j�A��WG����[�������(}|���)	���{='`��3����'��ɨ&/U䛷l���7^}�%�m۹KR�4xVצ�y��������.kX/���Տ>���ޞv��Č��x�V��ə���2���9-Ub���ӭ[Ŝ��+?�/���C�!������]�	�o���ja��KRzZ�����U��S���ډ��>��8
��h���3��͈M�Қ�ҲB��7bߞʍ�Z[��щ � y[rȘ�s�J�s�a�C[s5b�������7#=#[=<����W*�\�n�YbS�(�qQ�1j�rK� ���`tt5u��-��upv@wO���{�v�b	GdH=�e".&	Ǐ�VȻ�넁Q��à��K��&P�F3^�m�w��/�c�-jIQ��0�g����s!���C�QL���䈪F�0��3�{6m�O����׿��Uk�p��7��r��4,m����;�]q�-�(���9�����{��W�"�lm�cq�@)�88`�<���ŭ�̏��e�a�zIu��O#b��8�vj1��f�AWG�ʳeg�j<��~;{[\s�D.ZZڑ��
#���JJ\r�@WO����z�We��W$��s�A��* ���PVV��z���#��X�[_�++[�Bã���3�%����->s7�7nܠ�A6���ڰ~#lm�Q������Ρ��A�n�C\YY������Qd�f(�jl��4x||,��b���&p���	{��-�E�����BE�剄SI���N���F}}�1
g�M����9�!��5�?��c1#����m:>K�B����!���}�{�vJ��GeXJ�o޵��}�7��~�� )���z��y�Ԕ$[�͸9;H#��aQ(������3�ʱ�I����-�$zϼ��vfjZU!�X�Q��� .!F�:Xj�����a���锇�1��TVV�yL����`dԌ�%��w�y+:��q��g�X���=����Ț�����9�2��\/՘5�9��rAyI)疱v�F��y�����i�'�  4X��5�u��	��~��s�'ùr�<>+�q�YRǔ:gϞ�����.8�Ҿ���DE������on��ݻTᵶ5i�Rvv&|�=��ڤA[6��	x�r�*��Mt�}�    IDATb�[��I@���M���_:0$H!�8!�� Q@��6w3�y�����Px	��߹��4�Pp�<~���!0$TC4,�ã��Zp���];�ڹ9����瞻�����Z\L�=�����b!|�T��B�i@��P�^� A;� Y�%0T����K�;	�쌥�ƶ	~Q��"�o�������Å�|���	�lmk������r.{;g�Whobb,||=��X���J�'�a���hjl����d�����0!�C������������3ib9����%-�����(����qNt/`���Ԛ�[����b�r diyN}���q��Vi�#C�����0a��yV�6��@{�тr��Þ�;QTxA�CN���M���|�hi�c�X��RkK�e�U8t��E�c��˽XDM˰8�!��2�:'����ɿ�3��Sض}�
2>�>�(�"�T0�@�vYi�ٵk��ܽ{K�e녿�p�W=�FDX����;�f�m_�P���6=V�`��j&��~�Ӱh0�r,=+e�yCX�ѨX�34u��������
o�{&���U�)�-g�4l�U�p����k)�6_/w���T�{y�k����a��y�A���#�
��wȫ�#P!f�νpqrAW5��T9�����/ �DĶ�V-�U����y�J5Cz8��ҥ2Mtt�������	q	���vk�j[���/�������HKM�����VS��ø�Y���b_
�wVN�6���Iqn����k	s��FFFhW�T,,�(��is�W_~M���=�nz=�X4,z�'�|Rw�"�@�%�wV���sy�6�up��ˇ�_|��G~�B�|�051*q2���m�mnI�5:f�+���j���(��k�"`����s�v\������k�������n�I�U�55���Y�F7�1�E��s��'�=�����+噹�		�qq���k���X�ё��	Ji��)��������N�Nѧ�\��Cf�A#��a�<cc��y�:��cc�<����iJP����~^���Wc�#_�p!Ar��SK��r@��V��i�|jJ
��XnڰQ�O�C�)���k��9�ឞ^2���c��lx���K�^���朤/��YZ*���/wOTCj�%âX�a����O=���(����PH�b(<���֭;��w���W���������\��11:$��-��8�D��aXn^�2�֎vU@(i<��@�Ke�dh
b�5l.SZ�O~��,��)$�'a��]Agxsr���������	�����PK��z��i�������t���4��βn�z��ŕ%���RR�����.���
�~��'����k���KPvN*��!!p#/��s�X�����3Z��1>6�M���QZ�		��T$DM�z,,-���_������U,1�!m���na�D�#҉��Hg�^�E,���C��\~I�.C'�-<<ܵϚ8�-F���}/'��,>|�#�b�/�BF�K�Eh���GbJ*~��*j0�'�Ei�3��v�����{��]6�����v��w�����IÚ6�iI�����7���@o������^Y=-�o�o�I�/~ ~у�[1Y������1#����t�6o�(�z��� Unu�Հ咠WWO�ϭ���Ganf�7�W]��$��֭�5��^��#��jM��N���g�hia����>] ���E5t�
��֪=!%A�`�<3LS������j5?sp��ǎi(#!>s��(-)ן��6��R�}@iDRRRR3qFXP?�#��h���J����"ۂg����Ks�|������)B����3�������ó��QX	�w0�gضU�s`�F��=?4��gω�VZV��e(��а�(��PH�������A��)��[��_�(;p��߻r����֡C�6�{��︹8��`qnZ����P9����2,V�܄���B#�fK�1�=��� �O�HY�0�OMO(tw�Ԁ����V7�0�$���ǎ.q���xxyr��V6Zm��T_/��4��}�i�2�Ƚڽ{��i��7ܨ���O�.�D��ǀ�摖��q���"�vvsU��$߬E�S�R�b��̦VCdx0���no����T0��PYU���p��,YXK[��J]L�ɨY��AR^�4���y������}�fm{�`�̜lKL��rC8�ȑ���͖�+W���	���f $$��#�ّ��rx�ω�_�ޝ�%�[/�ҹ�;�|)�Io������Jo����۹�䲆u��������--������a�e%�L��VD�����������d�1��r"�އy��F�A�+N���W]q=:;zQ]A�aW��))��J���SŃjj�@sS�b~vv:JK���7�o��^()-:L�ӑ�A�'�$^FH�m���5X�GDG	S���u�e>)�t�\��*7G:���s!�)�̅����"ͫ��$y5�@���dgWg�`y��-=����9LLOa����,�χ��5r2���g��݁�[��9w�X�bL��`���\\UAK�/�{���O�:�_<�������h/o�vP��kw�Lf�eg����>׳�Pp^���׆������x�7pӭ�	y����YY�*����r��޵e��R֣�|���!���PX[{b�n�zY;M���h�&&'�53 ݂a�R($�"Q�ZFG���b��$��Ŋ=:�{��6oވ�@���DH�OHH�����AHx��T���ΟDX8���u��nW��z�8q�344V���]U���8v
�6HNɐ8~�(9	�Qpq���S����Wgxz����VJ1����5������Q��i�䏨q������f�t���?�ѱ��m@kW"c"����A�nMI�y�8ȽgۋMu�N���楼��UU̥.==�8i��%����5��L���lc�φ��$Ur�:C!����!io�ubXhX���>>_돽�ꫢ�|���`��2f�S����܊���7�~�y��=��XG����'�~����'9>Qp���e��C+��;�g=LF�&��*�c�1I͗�w'b�e�EA��\��	��Л?v�B�-�ܬ�UVV�.}tT�ɜ:�m3�>4�5^�����x8�Hw'���-p�ȗ 8t��7`��M��jo@TT\�e�]�XX�@pX,&��Z�9aGX�?�<051��s'q�5TU�����ظy�F�斖.2�1�W��`��tOO =8�K��t�����>pquWA069�؄HU��%g����Z#�FQa�
j��t����]�'�6�*Ӊ��h�E����L�=����hli��G��f�Fϳl���A<FN8�ϴ���Q9/�O y�Lk8s���^x^ľ��k׮��<s�f��05���-7^sCHH�!�u��!�~���|���Ǿ�N��W(d0�Ǣ1�_+�YXBOo?���eº��ζvVH�!uM�X�0�Bz�!	e%��ܵ�ҕ��Ğ�*�
�p;k;|��ocr|R\!�ҵk��߱!���;;��y)T46w`�<���dD�����}�m�L���UZ ��Ճа8�Z��O]@o��RR%�A^VWW�c#`cm/7�wv����vNHHJGcKںzE�c5�Q�q�����0�Jl���>1)�vN�(��DOo'�g�1�h��X���|�|��; <������2xD�KJ���� x�+*�u��xd�2T����)zb�`tv33�_N�L�6������B9/���<�}|͸�8������5���.s?�$�8�����.��m���۳�/kX������o���K>$�9;�J���ɮ�XZ���Ҋ��IMRrKQ|�G�����;?<o�%>~�ֶv}�D��&Ym��Q����Up �~���L���	cb3)�����
Í;{b��]hhhAQ�x�8!5)S�Ø�����(��������Pܔ�ON����
�}�X�.W"҇�[�֭;����:�u�����.�J���s����,m�(��|��z���KKK���0�M=��uENN�<PO��V�Qm��.��������0�`��X#�%����	������"���6�6z8yμ��q���C����7����)�%�aP��W�'�د~��<����;rWP}}#��Q\Z�~�?6�[�_�������{��_~��'|�����+�i���I�]����jw� Lc#pqs����Y���F����p��p	��ЅyR����a�	��bI��썙'���B�f���:�.joG\|���"mĺXJ��'!19���?Tp�ڹ]���M�ڀ������$4�u��4� 5s�����%��`��1!V~�^~��FQa9�m���)n�-U��ؼa��QVV���ARzU6�9������J�,��Օ�{UYTu8a��;ב8�ss
mG_���/�\L�I'������������&p,�x_�aS�~������XH]Z��ѺI~^oo��a�K��#����u�]*Њ�˴�������g��뮹�A�.
_���7�99���}?�sqt�����}>�5hX�mXZY��iT:��{�@�\D��@�F��_|H�Ľ8���P?s�� c�ǻҒS�Y tvvi�0,,\�7�%�w�bdӚ	��,�'�ٌ�� &7�!4$(������yvVTe~���$�{�p�UWbj��FeNz՜�VVv��$���:=/���"��{5�H��Ξ!ɑ�x9ٙB��{t	�������:~�		ؼc/��eؒ�����h��P�;iP4J��qE��1--ZhX�|�C�)�4�HV�N��1��Į|t��w�X�x�!Rf��E�2w��T<��s�\�����II7�h��[��έ[7�yY�w�c�~��iII�?��#����=�$���0/�"�K�kbrZ3fܳ���P&�A�t���՜��a�|I�#)9E��?c.������o?�L��W%^�؈����y�9��F����I)\Nl�Kyp߽���-((�@�={E��X:+�]۶�����
�+8��1+�6�#�wi�@4�1�q�6m�����$'�(��h-	{驢ɴ�5���n.��ҢX�d�z����; �}�46/�P�xaNoCڴ���E��H���͛����ji[P˝Mv���^	��5ɀզ��eC���Sސi>������l�)_�tӳx睷�{�9����c�)�LclΛw��smfZҗ��+\YY����?�ezr�/}��uEy9b"�&T�!"fi�eJsKKZ���ӧ<�^�����ݭ$�7�����h�47��$��d̷�[jcm ���q.q��Q
�/�0�I�i�hzLT4��je�������,"©����%j�b|�M���_��Q{~���
��b��eK����Phkkm�`723R�+�?����ƤyF9���DI����	1ѡ��1f���p��㘚_��E���Zc6@4j�(�����E��j�����N�ǵ�7��^��k���\���%�=*ϔ��gȞ�y5յB���X	��f���1ml]�~�����E�RW�L<p��v/Κ�cbb���W�+++�����"��~���l���_C&�ziD�Z.D����	`B�������>0`&�+�fX^�Z��0|@�8�b<�%�+������ػ{/֭[���z�kҙ4#,�p��U�{�#9!Y!����g�e�Ftv�*	�����5I|�8�e�]�Q��\�m��M���D_{7�*����
�<5#9$k[[��䚏�`Fh�?��Ŭ%nE��ݓ��㨩�N�>�2\;gi�k�3�7i��-��АL�gQXZ
7O/���08D�/c����g2Iy���k�
P���C��{~�S	��`cnsڐ'�)XZ�����_�Ԍ
�@��K��Gj6�92P6�����i�W��%ģ��]�Gg�p�fb��=�N��$$$|��;���~���Y,�޸�h����QUx�E�h��jq�G�)i�@u���I�b�E�P��%0�E,�FE#��������;]�d�6
����Au�uuje����������R�}l;�9���h6�[%���$P��c4���.�g$���}��i�ERB2B��5w�����p+��\%I/&*�3(.:,�#*"Lr}S'&g���p��9�;���Xx�����ь���&�o��
���a�07/H�9��ł�H7�^捬�l���h�5�k�+Z�{i 4&-x���z��P2vn3���iaq���ܜ��� ad�we�98,D�kR�;w}��o=��ݹ{�BNv��ݝ-o&&&v\6y���U^^���o��������)$��hM�̔Yo��g���/�.�����N�>��δ]�pl�0����f��0�d����SE�[���x�U�u�l�f���NN�%�9"���F���S+���{�,�w�BR��]��]|�p�ԗ�La�aZ��œ#�����~ >ge��0��~8�� .&>ޞ�;��!26Q\s�
���8(w4>AB���u>4dP�����=&��"�'�m��&��e&��c$`�����ǭ���[u��*����	��i�4*�g,�����#ՙ9$w�P=�z�4,z::b�T/|���{�^c���N2O4���^�4�˓���hoo�7//���_��}��ǿ�����KQ�y|��ad��)�$��P�K�Q�c�nJ/RQQU.D�����h��>X�r������A����k�����[�a貙3�ְ�<s�rv�i�U5@������Z2O�r�����6���a�����}���HCTD�d��:	�)HLN����0wkiiFKs�<8!nf��X���8�#c���vqM����j=4��Q�΂��;��Ƨ
��L��t$G�x>��4���B���c9�C��qx�}X4�@�ת�9*����V$��_�0J'llWpe��eoO�v^t����`9�z��	�q��YS33���Ru�/,��䬄H�F�Z��Z���=G.뱞y�;~����x�w�x����y	1Ѱ�������L^44E]�ܰKLLM���\�I;�<��n�A?�0]�1PY�C�m���0��m[���� *��-�ʑ7����w���q�6z7޴۷JV���J��l�>zT:�yY�hmnąsg�� XY.���#�6�T%&�����E���_��r:�ʎ��y�X�
�f�*?�/�;;���\�����r*���4iȄ�I�i�f��A��#&����hnl��j|l����)����T��a��U,�3b����X5�����-[7�(�l��3���/7[5,>��C�+���czj��:z���@Ҝ���2��o��54����.��� 08D4��¾�޾{n��w.kX�}�������
v���ƃ�'[[x��薲�X�[�'�a���8{0)�,��TΝs7M�3"�(JVA�0���������������u�Qg�UTL��b@ń�HMwӉΩr��;w=MɈ�w}��%�T=�<���O��s��"QM� fa+���w��Zx(��s���/w+�4�ܬR��SrVd�I8��ذa�J����Z%�,rjT�P���Ϫا���;���W'eA�E]b���?��s��Q9h�>xP��-���'�Y�~�,X�H�>��ڽ_���g�Ҡ���_ʎ/����l�_Ƶ�"19z�V�5��V�:/�7-M�
g�'4��p�I���nڱ�q��͗���n��@̈C�݈��G����M,��U��5�k���j���f}��gN5`2��T�s _[�Nׇú~����š���O���Q�G*_�`��oi�*M�{��Y���믽Ҙ���Z����N	����˒??�����T������jٵ�̅�ъ(SU���Bz�!�g�-�D��*3eDN��?X��T�����v<B�ǃp4�2�    IDAT��g�ƌ�ׂP�	��-^|��w�a�HT큒�|���[�d��j����[*IK�eP�`�`?v��h��[�J1��"��e7��AUP���83�%�fƌ��ߞ��>�_Ǝ�(ë�+h���+CG����Ƹh��O�3��t�Cw����R*�Tj+G*�	���p����R;�QQ��b�x������2��lٹ{�:-H�M￫��ر�+�Ե�*s�M�`�,V��C>�c�!C
h���9��tV�n��<�`C����ސ��ٹ{���5�mw|G��ˊ�O-+.��u�-~����}�]�l����������;�z�Q)/.����BR��k�-�@([āwH�F=�ťf�;�lX8mDF=b
Y�G��������D���fj���/�T�lۢ�� (���jV�M��v�Q�j���H���m��њ:ٲm�J��G�7���'�-��+�u��|�^οp��rK���Y#ݥ%嚲����Cd��3��X��R�֩��y�(��~`RN>c��(��G�u�3 !�Q�FT����aLHT�+�uR�]���F*�]��:@b��� Y~��?�7o�����s�IWG� �B�^>��̞���]�+!�m�	~P�4=�5s����{�g���
U����=����7���R�������^V,}����g�u͒�^;%��������V<p {�E��K/�_���X^�~`q�~_HB9XI������|n5��<�'�^K��8q]��*�裀M����������N���d�K=��`�2স���Cn��v�	e�/���o����wɎ];�s���EM��֒���R�/(�76}���O�A8��4(���4��7��T#�HtcT�@��_+�EL�F� Z?�=7�P�I��4_F�������|�[�$H��T�h,��뽿�C6 �f��c{�ٳK�9�l@����� �z�v�@����O���?�p�s��q����'i���/w�8��#�\���� �����/�+_&����������M�\�����ߗ_��ҧ����ˎǢ�_�#�~�����2a�(�S>o���p\;�9\��5%^����������U��-Gd��	Qy���Sj�h�?�X�8�Ʒ�V���.q,N���W�46�����پu����x亨��,��"��Ig:*�Q��E���~6�K��s���B�u�S������q��W�<ҭ /G�Hs:���c��������$+ �\6�'"���m�a�O�f�.�W�M�����t���g���ix��;5�R�f53=ph��`?~����~���ɓO>��U\:H<�l9��	2y�H-�}����x[��0Ϛz�447��77HYq�Nwݵ�Z~�O?�!cF˃?.�mڼ������W_��)�u��W�}j��/��������JN;\~������C�����_:;{�sN���JVn�J��L�jy��� ��ۥ��K�3��֚�[��|��#�L� �9��/���d�mZ��L�B2���TV&�.�Tv�?(k׭S)�a��M��L��s����Ͱ���ɰ)���� a�x�9�D���TIEJ�(:����HI9\�:��E���ä��A�ؾE�c;�4���-M���իv#��ِ���\�M= oyy�L;w��_'5�����b��(�ۈD3���~Og��ɍo��a�i�o��G��*� zy���(��xJ�l�p�3g��|Im;��{�G��˯�Ire��4��u9�G���#��]�����'�?�U�n���n��N	�?���~~��������d�J��}O�z�!9VsX�"�hB+Db	�X<�Ã(��a�+�S��y�D�l�d�9��-Ǜu���;o��#�?j��������dsbtntC}:��S�����ԛa�����:ݜ���+vT�T�dD���I8��͛?P[b��!�z)e����x�t��HmM�0��y�ހ��{��qcFK~n�7�i����H_uf��\)E �5�Eȭ2��pu���(���=w�I�BRq�<��ݍ�h!/�ENi]���DJa[YE�H%԰�����D�c|��ꨜ6�L:�J��,}�Q��k����/�2z$=l�C���k��˭w|G�͞'k7n����@�9|�5W�|�ճ�?����'�X���u�h��S��w��-!����r���U�b��wH�^N5 M�}�445���B���Ԗ@j�JG�+]@�z�{v��@;kH!dʏH4l�P��$��&)z��y�w���Bf��Dx<>Ge��5<2(�B}�8&�����X��&_c7�zH�]!&����.bɨ�A�$\ow�JF6�z=BP`����d��~�i�ޑb}򩄲��.T#�^XR��'{�}���nBZaRl~�C��1cTC�9R��f�8dH<��[+V��k����ث��B�s���ʒ��G�����~�~�k���т�C��Ȳ'�p<&?����;�HY��·E?|õ�v��O�
�{d�E�V�Y][�T^u_�L3Ln��
�����ǥ�}�,���^5�.�����wu�)àD��>p��bhXox�
'k�	j�a#�
����nj2����ëaqh���jk�ʤ	5ZNc~�&�xG���4#=���ڮ� 2C5��ۥ,�d<���xr�_;��'.�=c/*�)+�5mz���њZ�M�`0�ic5������oL{%޷[�^$��0_�����5��r�����!��͟�k��+�����A�'B (AO�_^���}����r�d劧噧W�W^"���5����.u�}�a��+�o}G�m�D�xv�D�48��}�U�r땳N]Wx��+<���g�Z�lB"�/�u���o��W_xF*+*ts9���a4�Rn��F��2pQu�x��/���:���l-��P%�����3�A$�EeH7`�o��3&�92�)� TA\��raT��>4z�3 �Dl��fO>���Ch�{��qzm��hB�%������\UK8|'�Y�0���;N��ﰻx~���z��=*��8ޢ�5�f0|��'
 &	�����s�齟=����]����=�� ���|�r=Կ���5�⠣����MP� ���~���o��:9}�ir�X�|�m��k�4�����[P([�F6m��T�%>{������;��y�\!�zl��g��;�4B��R��P#W]z�̝>U�z�AID��(?W_+�.�����s�t��̢ v��P���}�YZ�k�2l6�����\��f��x-/ה*�+���R�-��4+�0�7���n��wޮ�$�$�~$�Yxzp-�*@ӱ`�w�������/0�s�H�vs����ڝN*���C�| ��9 ��0�f��C��#u ���6pϰ�C�5Ƴ3Y�*rz�����.֘�`�����[����A���J"�'�?�F{|�\r��r�-7*#b+A\��Ͳl�
Yr�Mr�o�u�~.�=���G���i�q��o��峷�:�����\�ܳ�[��T�8$&�v��'?�c��u/���R���f�n_$���7e��MMz������P���؆ @�1:27��kz�J* �J`�8�����2��5��J7����B��CGnik������C���x�R@L_vz��N=�LI����W�� %p*P��P��H�@m���B7�#�l
f�t����O��Gꚼ�8#�d4� ��W`B�v���%�/����v� j�y3t-�ǰM�`�EG�r�4K�`r=�����Xحعm�[���=$[�~)?���eA�ڣ�嶭R\T +�.ӂۻ~�/R>l����*yi�f�JL��pێ���뷯��������V-Z�|�3G�Z�v�i&������a�}�r���ʣ�Yzښ�% hP]�}}�?�O'c��)f�Y $���>}0ʥX`#\�	���SC��j�#�xE�q�㼟I��)���,�O~��y�۳W�ƍפ���t���s��k�F���j7bS�V����Ca#�D���D%���|�Mj�Ca3�Ν��*
7��x��\(�&GJ���!���Tx�֭Sﶼ�L�˰oR�����eݐT ���5�q��\��N ����x��T>w�p�NSݺ�K��{� ���P�e�&(˞|B���Z�f�m��ǻ�O��=5-2h�Dmz,]�v�pɜ�p��o �#+._��ŕu�Z}6�O�M��.�p���5�O~�IF��UKe԰!Z-B7�(�"qc0:�J,!�L�p%���� �H ��< ����,v xl��h�~�'���c�Ш%h6�?����WTh��\����ͣ�ߢq���5idB۲��?_#�RT���P#�`$U��1-�`)���3a���M�D�?��#9z�F�tt��O�)��{瞐P�	.3l|�nh��A�Pm�axc�B�/��P�XX���X�<H�!�h=�` 4�1��z�y|.;/O�RR��s�e��e�5�JWOT�o�!�W�/{B���������O[!Ͽ�Y<�%,(�X�Gl}ͻo�|�w-���)%֟Zv�ҧ_Z�����W�P8�1v�=�[Ι2Q�w�yf�����$�:��]��6��dJOdQI��W$�i�p�C��Ԑܺu��g�9U�dMc�-�Dܳ�V�&��}�Y0b94�3�B_������/�S�H]N��Ӧ����rO�0+��b\R8�H��w���:G�{İ!����ݥ�h(ϴ����מV�Bx2��暈@��A�P�m�o�n΢JO��\�m�����%fu��EG�B#���P
���A`���z	HP��8R��	�� ᯑ��@:�UVʄ�N�a�%��7��nYr�2d����&	��e��=
�[n�Q���6ٰi����O����/*�P@\���zv�p��[~�dީ������,z��c-����+�}/E��d�[��~�V=�B�^���^�ɧYE���b1�̉�3N��!b��>~�X=5~���g�y3�U%���_0X<T��-�CҒ�J��&�b#�F���Q�%��4�S���K�
�����k�r���7�=Z��Ŵ�K�!ZYw;$'�Ic��Ї��,H��@����D�y�ŒL�ڂ���&����cP($9����E�� ���:�L���J"İ(x:\%2�LP��F *Nv�>�yy�}��SQY��ֽ�a�D򃻾/�'M������/�e7m���w����m����U>��F\�RI�=RP�/^gL����o�t�?���T�ߖ/^��e��
�uШ7[B�����'�Y�"�?�@>|���h�+3m��͔z
$��G���A�c�(�=Z��K�b��ӕ�	0����M1 �#��<L����Q���Rs��j�p}�l��iW� �^�@�Lmln��3gi�!����VAt.�J���g�A�>���z3Νn<R�_**��j�P-.���ƖF��:i�Ʉ�Hu�za�J
�.<6��b�3Yv��󥱱Im*��I��>ߢ�9|��b�Ғg�b���d�vܣ�>�������$� � k^\V��T���,�X��Ѝ������d��?��Oe��)�����?+��v�+*��Cʋ$ng�}׍�͹��]�唪𯏬��U/��i�T�K#���R�>����x�\0���M�ɪeOJs�����ޥ L�L�5�,$eL��<��Q�8\��}�T]H�ˡ��_��܌��A�ۨBN��gL�ů9|X�C ��� 㶼�T��	G
VUUJ�y��h�ТU��S%S6�T\9D�J *�TU�|'����F��ʖd��!�*���Q���u�٪�yNT���ςT#�C׻��f�� �q=t谁�a%E�j����ʕ(ܡ�jj�FH�R�����bWaR�`=8��۔�6��w߭Z%ަ���_�R�@��˗�4����ʶ=G����|q������)V-T c%���^{�������>:%�|��EO�z�����8�bwy���IgW+cV%�LI���t�ʯ����]6Y��U�x]:%�����5�%����8�Yغ�G�$c�1Bk�ּ��ģ=�S&O����ba !����X��j
��u�@KS�*�����U�k�;��5���ϷnQ�S��i�d U*;��]����]&M:]�T;s�I�0���vf����1z�hٵc�N碷D �'ͭ����A��r�7C�x��!�:���3a{Dզ��}��� `2�5R*}�yN�����$��T�\l��yV�P9D�@0!�~T ������'v�GhŬ���ԖL�vT�>��Cړ�NɹE�r�o�"��~(�`�Dl>�C�����+!�����_9��_ѩ�Џ,}�G�=����)�r�لx~p�
�s$�u�ϖ�(|��K~��*;wl���xJڇIL2���'ݚ����xJ�����Po�t�S�����O4�3w�l�q��������?���k�0|n%�Hs�O�P&&�m�:0I�D1�����| ��揶({󒅗(���eC��G��w�R)���xR��Hv��	gd�h��F-xE2�����v}v ��@��TRPUAQ��ܽk�^��16�3	�^�g�`�q2^�����Ŧ��������� 1�C�2ٞ��!>���Â^\f�F�P�@C|��vG�9g����{����4�9D�J%j3�h[*!%Y��NE%�w���Wξ��Kn:��zdٳ�Y��s��6�RΠ���$�j*'DV?�����l�	c���fɶ�>V���w�mC\H]|zl%��aʙ�5�%��uqP7� ��z�����g���0�k6��Y����4����E��A��4��	l�����u⤉�) a0����B
��.�[{#P�Eo�
([&A]�Ą��	���Eer���$77O6����w˄�ƫ�fz��>�fNs� � 0� �0@B7>$6��<�@���L,.�t�H��F����_���l*_�/�^}M������!Cu�2�z��%+�|RUfy� ���7�<Dbɸ�k$=}��]|�|�KKgX����)��6�-�X�����mX�^���=�-�DסkN���oZ`8���W�c=��3�}����m	%���l��)g��*|���xD"=�i�k.�'�F��;w�a#��c �`XMz:�<�]Na3�į����o�Ǆj\V�"�g����"P�b3
�l �gn?@g2���ڥ�2�����F�#�f�Q�oܸAΘ2Y�3 `�.����k*��@'�S�ZPP,=}��t6b����F�=�;jҤ�D=���f�V��}r�++�c����᰸<.����Bm��}��.|.\t��s�=�ﯬ}UmC�4g���~@U���*��{�J����C9gڹ�	K_����������6\���.IgP���S��ʗĝW)�P�DRnI��L���uIq^���=b��U_{��;~����
�y���_���k�g%l~�3�	��EE*Z�����n;&!�Ȓk��`��e�4��a�@��A}�1��,X,�9sgɬ93�ȥ�'���+�b���D],�� s`F��T� ���6 adZO�n��O ���7���3�N��<T��XU�0��xLب�\AZ���X�]��q&�9.����&���9I� 8 : ���š�Ə��΋��Y�@�?�,��[���P�H繐T�� �E��;��h>CD��8 88%��z��$��y�՗�����v��h����(׊�]wO��y�y�N��g����׼)O>�l�sX�y���)���B�����W*"n9|͢Yw���o�Rb=�l����~���G[r �F�]�;͌g�-�)���z%�I��C2��X��r�$���}�'b��Rk��%��&]<4ꢵ�U�#=2r�p���d̨qj���� 	�t9�z�jA� .��D������!MöF-����č��ơ���ͷt� �%<�ʪ!��.�Gl[H�    IDAT�����MF� u����Z���n�H*�4�l�p���P�Vq�iދ�B�qM6)?��r`��>��{��F��Ǧ�9�����x��b?� G@���s%F7P�\<^����/��a`'�#��l���<p�_t�o�q�\y�b�oJ�Y���}�E�"���O����d��e��eoM�Է�K��^��Ej?k��C�Cq�#"�͇�_8�Οܲh�)��t����b͋{�4e��xb����h3��Q�ϧ��X_��q�][2N:m�\�h�47T��m[�edoW���wTB�sLYRK[�tt�K,n6y�U�*���CE5�����W���'5�B�m
b]^}�H�_��J�TJ	~yyf�6͵w�Ϩ+N>�&�ŒI�7n�p�$�F�L> j tU�lI���SA4�5�w�<V/*T-/��{U���p^�h%������>K$��u9\�
����?��I����P�����U��	m�g�c���x�\uՕ*�l6�z�{���7� �}f��|����P�j�_���r��C�<�}�N����b鏚��8Ln��b��?r�%��������zy�C+V��Sݜ��~��"aq�l&IOj�s�]�ݔ]^��뒮�c2m�D�;�lii<"�jk�s�=*�Sb�= ���7�	�_����0Q�NDʉ!Y�m�W׾�j��4b����t�p�yPB�H�W9q'@�jD ,>�`�'L����:)K;j��OS7�bT�J��kjTHC�� ��B�`/r���y� :D4�r�Г����But ��ye��.�=�ZV�|F�N�BP�ĵ��	�}ҁ';=�/E��}qydŪ�ZiCWū��Rn����`&<�n�X����2*Ə'w�s��r��g��OV���%9�c�!�����W�}��X,Z��P������.�q��z����W�ya��c�1g@����]5�5�p*MƖ�K�m�d4"�xJ�%�=���(�'��E�Jw�qٷ{�><�m<&bs����Z0b��x�V/s"I!%���P�l�E�	�D��(��5��;�g3�@+4@Kj6� ���b�ϛ�F�
����I�iՐ���'(���%@CM��>t�I��j%:4Ж��qX�oX/@H��{@�����>~�L�	ܿU�E|kժU�w����a�"��G�1�(Ɉ��U�B9����������~_C:H�H<�=>�l��[�A'Y�,u���Ī5����Q�RZ5Z�	�=�$6�����Q��s��ў��m8�d��;�XO.q�cϾ�fס�܈ݧ�����,�Τx<���#a����>q�D�{Z���I�_0C��y�D�:���!Md9rT�Ѹ��sL���S���ր��ף�b1��	F+F ��ުq ��JD����L���z,��\$��T��1S ��.Qu�K��Y�+)3��h�ҟ'��$`�Ѻ�oHn��5$�{0��L�AYCg�*�I7���I���ܗ]AJ��J1�҉�� h��Ͻ^�>1*�x��D,)��'�-���?��.��] K��VG��u�䝷7�;�}�3�n��6�����w�w��Wٱ�F*�M�a�	�ʎ�{��Ϫf�n�L�[�	I�t��.�x��z�%o�Rb-��Y-q͞��*�h�ʰGR:�EIu .�ww*&���A������}NIFz����̜6E.�+Ǜ���i\}�:��Rj�kh�S���4 
� �asi����5�B\	�X��fD�Y��B��d�s�DD@�D��b���63-É���Tĵ�7���Z��I k���˪_��J9��9 �������Pz��Bb�q-��F��Pf �
m�2V�*�&���l4�Ζ��V�`������r��]{��� ���խS-����5r������@�����_�M}.���P�I�d�`~�8=9x�*ps�h�s�緻9��v�%�YW{ݢ��������za��漸� �_lɄ�I0�$����|�TL;�66?7;G�a�DL�?�p��9y�\|�ij�{�J�c�,0�j���tjŪ��^é�C�DZ0�6�`�7�d���Qj�U�50�2P[,8ҭƬ�I�l<Hy�G��� �8(�!���ݥm {Lal6�-/?WZ����_K)C�!�;�����&ث��sm6�<���W�O}�DVU�-�F
 ��g����u�vN��{B:!���ە���֪���Wd���d��g�-��)�ǌ��ol�ǖ�������W��$;�B��,�-(�]�9ђXXY�f�r�x�qIt��^�p�w��Z�ꕙ_���?X7�U��hX�I����zl���v5�����*�x�\�E{�O�	��͒��h�XX;�y\&}A�&K2a���W\y�2Nu�oc���N�."���	q�q�� N=j��e>��)��hHQrp��0z�0�9�c��؅ �HTS��J�ˎ��(�M��~�Cage~-�gY���w
'�3�0�6�����p��OLC1.�O�����a��r�`��[�h�|�����%}��:�q�]����i��)gM�o�C*��3�o��V>'j[d�03����EU`a� ����{�A�n��̞0����n��n޹��۝�`�/z��W���U�*DbY����C�8ER1XtF�љ���[)%��H,�#�!�t��K_o�L;{�̝}�J���>�V<�}9}~��/m&�
�����J��H���k����릱�D�X�7l<-�_�D^��G#N;��X[_��:�@t�wj�ic�Y�l�Ƌ
M���n7�N� ,�ʱ`�֒�C����	��,�aAU��˖~�^K)�,*6
P�����V���U�6��h9Dʍ�����j�~�m�̘9Wn��{�	ɪ��˪g_�#�M�/�J��3ck���bP�Rc�7��P��������j����n��|3�V�~��V>�җ�0�}�P�H,Kf+�X�M|N��"G���a3T�+&͍5RZ�+K�[,�F��c�u�a��RG�&��s����Q9l��z�n����`U2א&���f�7"Qo������a��c{!8yxzx�4��R���+�H����#}�I�sF���稤��s0�&a`�?ܫS?|X[4�R��p�)��(5�il�mFc�!� ۡr��Zp��`�o���������O����,]�T���-W_�Dn��M9d�3�Ȫ5/K�|Y����;��"�8(����2%�r��l:;����mW���%���p��so���Kן�x���~h�/��__l����W�d3fΙ�@+az�lI�S�,&����mw+����M��4�.�gL�k��ؽ�0K9�H��� ��7l&B�H�Έ��t���93��r�������rE���!��6c���2�T��I�.2:���D�1H%����W�54�.���d�^#�P!Q4=��k*�`�СU��A���mmQ:2�R�5�^�	�P�	���5LZT&���>���5m���ET��fLY��5u�+�����v��������)G�{�_�^�(MaqQq�Hjڮ��L�ZZ���Q)J#p�JT��i"n��a����qD%���p�g���߹��;�N��)������g���L���J��u:�b�|.��wIO���r���K��E|
�a�C"c�{�M�V�r��SƁ�=��ب�و�#��/P�B ����D�谨���FH6�{�E��o	i�P͜��A���0q�O�~�sO�*&�Cr (��������Ś�cb^��cb
P��!�|�6��� �4�G�G1�e�_"n�՘x�n�>\-k_Y+���N�_r�r�e���fy�����E��u�$�_*�LI�exU�4��H;�d�.�<X���>"1q�7+_R�er�n��fy�Ci`WS�U�s�7k���>�����<p�Ĥt�*��.�h��ˉX������;-!'a��,bW�S��5vJn�-�H�,둂�l���Er��)��gr;�Ӭ�(�y�'캙�
�S�T$i��Ѫ�@$ �0�?g�1Y���%�L(� ҂M�� #uƐ���7ޡ��@2�X��gΗƒ�Y�3��(�5�	��Xh���2��A���� �N�L{�y)�%�����@���TS �ռ������J(o���J\c��r���Hհ������G����ݛ+���s�'�T*�Ӗ�ʒb��n���CR���>ʕ=I��Q`ٜN�����)�A�x�Q��o�₳o��[���?��/m�����^�}����|��TH��$��k��n���N���H@r0F�#�pO�$"bû���.{BR�>	�"�ԳΑ�����@uu4��\�
D�!�1ǆy1��=j@��!��e����ץ�k �*�1b�Έ�9�KQs������Pq���$����B��s4-���G�-��Dc��:3<i����G�~�\�kX��lR��-j��p�|�c�@����M��7;��	�C}f�Br�{I�\��Z9���R�
���rp�!�h����K�%�o�I�/�T"I����3y��g��3)��6�����H�a�!�L��R�O߲�r��N�s$��@gU��h�.��<-���ݦ#\�^�${�.�{���|�W����g=���/�=�TjsfI���!��L�%�(*��ƈ0���żQ�^�X&�/5]�>�no~v:���H6�M���/�%3fM��B|���?Z'��1q���Ն�H��p��I�z����յF��� Os#�
�A����1�L5�G���&��-�����] 	)B�A~g5� T�;�����v���4����D1@��c���۷ɡC�ڱ���UR���U[r;�*Q9x|g�{���ML{i�G�K�a'l���=Sn��67�4�m<.+�{Uּ���̘d�|bw�%I���6��v��#	))�סZ8:99��O7@�W��J<i�`,T�j&;qB��$���p�g�t��.;u��ߘ��cO�����L�`%����Բqu[JR)6 �j��� �\�HI*[2"�h��b�����O"�FND%���\�I�&��Ek�����6}�y>��a�FQ}@�ZvZ[������6��a'�A��&�����S��\0����gS;	�D�����輑vx��5@m"���h�?o��!�*҆'��g�c�\@�{�(��^�%e����9ZA�TۡGi�tL^|a��z�i���o}[�̝'��|�������o,��"�$<b�Vv%�ɖ�X;����oV"e�@v�)��ln�l�ԛ���̫'?���W�T7���I9	RysX�c X�����
t*R>�Q2W���U���)���ɭ�=�������=���x��WaĨQ��aa�:ڕS������*'+����l�"�Ƅn�c�b{�e���xJ��C����!}�=��0��f֌�Ĕ������ !U���Ҍ	��ܢN A�B ��rl4��Dp1ǌ�> �E� ���2a�D=\D�Q�<Fvc}�l��Y�b��\r��r�e�ʸIS���S^^�Q��|EZz$�`�$>鏦�1��������TCYSu ���p@beg�h8:6"� ��8���"�rBY*� �Uκ�S:�׽1�/?�Y���P K�x$V2�	˶bQ#H-f��6�N���!�A���ۑ���6IƠ��HNЧ���5��ڡ������gL/S&MZW�9����z�MU)y���gkgAKR լ&�4���d��T��C��Qa�=�j��@-RH�a� ������K��S#�H15���<���ڌ�a�d. C26+L�\k�|���"���yc������u0�lI�;F!�<��k�a�G�sw�tv�O~�D�.�Q�M��!C8�b�(�T��HD|42).��v���	�bȦ���GU"� �qK ����U��|�mߠ
��zuOuS�wqzT(��- �����R�f�*��";`?�F"�vQ�*�� �)�A';%�IF�\v��=��m�/w�?G�	6�C���A�:HƎ*S�L[<)��[+����54Hck�3�@C�p�
�B$��	H�����Ԟ쀂��RC�B�	��!�^ka@�D9�Hk�!�s
<��|j�+m��th!��;T���E��u�<j���~E���U�k��ٯ�����BW
L���%�ׯ��v�������p��O9�F�A*"`Z0@��N��xL�ɨT�j�`�줁EKPKf+��:v傳�X+׽1顿?�v���rX)�I<�`ـ?�o�`��E�3ŋ�O&b�t���r�m�HŤ0/d����R\�/Y0"�ڕ�z�Գ�H]����f����	��?לWaaPrBn���*0ǌ)ϟ'١���z����F��<��0$�u�	��6��J6��PfL��k��kU�	c�C�gޯR'��3-�jN/j��l�����=����S*�QozI���d�N�KG{�|��]y��u�e�VT9D���69k�y�	����e)lݽWvTWK~q�$SH͐��̨N�?��H�0p��ƛK�{M�a���ⴥ��|kh��	���:`Q�i�_u�Y����o`7X�R��cz9���8R,4�2j�fg�1��D56��|L\v�e���&	�2��T쩨�#�2j�P�()Բ#��'CF��϶�_�(��G�
J�?�&�;׊ʰ��R�������UCd�Գd��J���Vban�ˌ ����H�S��ڱl:i"��@���K�-���#��<�tT�2�0q��Dy�86�0Xt�����P���̂|Uo�.Qu���:����KOg�Nz}���������O��.gO�.�8S-���7��/�ǎK��_N��<�l���@dI,�����T��Tާ��Rn��<�F�:���PU!��һ���++�+T��i����W�x�Sn��w������ޜ�ГO��{�q���x?�T���J*I� "�*��48
��&�e#�{2&��6;|�\&�D������|�c��T�²*5<��`�x���顆�@	O�{�$�҉�#����A�ԫ쏴ɘ�C5-O�jж��-Z�p�p�v~Ab`�0��0Ae�C�+[�i�r�a�(5�N����K2�F�E�K�\��yp� 2�>��J��ɪ�A���Oqi�aY�-1*�_��;��#^�sΓ1c'��W��.on�H֬{K��4�?�H|�\�%ą���1B6j��CZ#L�Φ�bL�8Rqq����(GQѺ��X_H�NS�	(w�*�Ƣst����ۛ.�y�-����oH�}o�_[�n���!b��gh�DhQ� Ko�N! �8�f�&�j��HF'%���?r�,Zx���*���-YA��ؤ�;,��|[6��Yz�6�-,v�_z�a�~c�;1IE�$��%p�s�YRQ6HJ
s�	����a:ǂ��*���=;�T�;���--�?��׬�l��h|C�0>	���key�C�]�	ɿ��b�[������ei���!UR5�R���n<39ɤklԁ�n٢�r����7A�k��i���c�·��g�wʗ��J�(xN���|/�k
�Ӂk4��ݦ�8Mi�M�8�G��V��#�g�_ʊ���	,�78 ,_(�|NM
e�(���H[��3'��_?���#Oּ����Z�nۮ��vg���`a��^���O�I���`&�`~2R+.NIH��ޮV��vȠ�|�}��2u�$q:D����O?�w?�"��S�9E"i�ݮ+��hQ��&��$H$���_�z;���/����&LT����&.4j�p<�R_�A��;�����9��x%t@���D���,��V����7r�h-ٯ�����b���p:�"���v�]{��A�u�t����O��=�KJ+$��KM]�lݹ[>���r�Ai˟��铄zz.� *�JHc�#��=}�R�`K�_R��%���@�e�d�W���h���
� )� ���T_[��3&�����[wBİeˆ    IDAT����^~g��{�{lݎ}�#�l�U$S��M`ɥ�YC���*y� _�V�yY~��j���j���P�G����S������H<�ӗ��qMz���MX��dB7��E_w����T1ӵ�qhh&���&̔X����Ə3P�UR�'��rhX�f��=���g���֧h:	��II�(ǞC�0^�O��(���,�uoO��V��C�k[%ʰ �Y�x�]�<������ʓJ8��y���DisI�Fx.�V��Y�Yz��y͡'D�Pi Z�F@L���d@��E���X��xJ����:x�H,�ǩ��ݐ�kkY8}�m���kO	��7�3����X��H�P$����&5����=eT�,�d[5�RތZ�+�\�&I�=Ӣ���Nm�&v������giu.R
Y���@�nI_$�iZ
m��X�ˢ�^��ߜ�u��,�0~�L9}���1��<!�p&U 6S4�3�V��qd��v���S���������>q��n�*�tTKO��낉��𑣍���&@[�9Z/ﾷY����;��
J����'_P����	^�`���0v��:Y6�gx�x�L�¼R" K� ���y/T������X�XRB�yy�Z`���?c����ђu6��4�3Q�~�c���J�".���4�H@��q�sBH�ؓ&1���)I�5�CP.��8�bT���ƻ���	
�fw�E���ѨƈB�^I�H�4�����%ĆS���aS��Z,�AR�HX��>-���� .)*�!�+e��Q:gO�?.�dy=:
�~Gw��tuIg��E-��so�{���>���f�$��qh$���Pţ���2�oϾCr��N�Z�x{�4�v�ǟD���aX�˫�.�$Q��X¦ײ���s�9��׏�N�n�a�a�-�
�����"�{4&���F���,$��p4��B��-LX�0�s����o��膵��Y7p�*LK,V4�VU�kiĪ�Z�J		W��Ї&��T#9�nm:�Æ �_�;$�c�T��C�p�&	��s"��ax:l�$��Hh�Kg���oӾX��p��$��٦��=��p?ܬ�E���KQn@
򲥼�L�����h{"�)��*qQ��g�{l��9]�C��@�V�HT	v���#����)��;Tݹ\��T�(u�CI����1�
������Hݘ���������ߕ!(�BR�L {at�J�	�B�qF#R�����]�*$	m�{%���b�a6Xƻߝ�xwKۼs'�>�����ŋMR5���?�~��Q~`���umU�Q&{e�*Ԡ{:@��(���s����IXF�%��%���	 ���D��a���}�C���Ρ��$,�DZjٓbw.S+�Jz�����v� �Nq��VYH$�pz���\��X��e֜v@��_\��C_
#��
�A%s�<��E��Qǵ�I%/�$�jw���ZW�T�jT<a�$�n0�!-�q�tk�A�t��f5��%^�!6ޠ�+�5���
�tĀ&I��P��Jqt��b0����G��<��v����fӖV�Mb���O�s�䊗gϞ�Z`�Y��������]�ǆ�7����E�2ExP<�#V����J~���jԛx�1���Ŝ�c3�9�0�|$$�K�c�$����4��6�8�nm�_+��cN;� HpֵYLT���ŋ�xIRa�r�ʔ4wk$��'Jʌ�nrq*�sڞ�sМ*�m̺�k��P��]&���PV�H���kݬ��@���FH��>��8Y� k���fTaTJ����0�b���e�*�؈�Q`�+�=�P�/WJ�Ms��������q��w��zy�������n�y���������x�e�7T����j;q��+}��x����$5i�l g����H���06�FKIT�d� n�y`8`� !�	�z���ď�� ��O&����Mɀʁ����N�O�)d�I�E���%�F�X�R�A�j�֊g�5���g$�@��l"���� �Ҕ����@X�_l� 7!�XXJ
Xx�:�� _�,9z����X��Z$�+%��Ǝ9g��ιæ��x�)���������vlޯ�Oܜ�4���dK�I�d]̴�����\�g��-��-�3mc�.�F�M�J-���CJ%�j-7����^	G�����-8鑸C9�Mg��n�5r�Qit�J5�S7�� ���YUNZ��1H�k�]:�k(<F�'���J��iڶ���y]���en�T�*�	P�z[� Z��8��R�ﳮ���L�
��EJ+7?OG3���p<9`��Ċv5t̞:���'��`��=�d���;U�{�S�w���&�&�n�8�,*�M��9��/=�i�nk�s��ǁc�ڌ0dQ��`��>�G��� ���Ӧ�f�^7+����[m���4��8Z��]}a&ZR�{�}N'Ϲ'(;ܫ234�n6�����l��8��#i�%�d�9Z��E��em*��5�t}@�{@�q���e�κ�~.C���Oڋ�{�*�Ӛ�$� �pi/$%`5G�X4�Qj�l�>+��t�3u�.�:��ٳg�Ҫ���q����<�tö=��)H Kl	l���k��ƫ VZm������W��c� �Y4����@��:3� 
L	zC��.+͗��|����p�C�ص_�#)�/�����ġ�:\��r&N�ٌ
�X�RnOH,�g���)�,Uh]G�Gz�^epچ�T�Z!+H�!��i�c���� ��h��,�e�uNH���T�N?3 <���cL��p���v��V$n�XN�^IU�������#���:s�?�7s���Ӧ�-���`k�����ﮙu���;4�U��a!�d`Y�&X�����<�e��V0'7}�-ᗄQ���Y^�$���S�k���*tқ�X����ʕC�M���Hg8)��R-�A�
'�h��8
��԰��d:��8+�c�>��=2X�z��*���f#͡���L�F�$�J���e~F�e8�6j��5�܉ ��߫�F�cE�`H"f�e�hm��c
,z�Z�,::ƺ��O��N��|Ѣ)��}��Z�iK��=�~۞��X �����X_U�'$��_�<=��Y`�v�?]+<��?G �R)�b����T�#�A��Sa����K_Aa�T�#%��˳�l��oo���QK�%�kU&����N��m�rj'$�ٴn�u,pd�[�O�$`��Ƴ@�A�W�w��9�j����!�fX$'K7#MӇ7FmJiQ� ��
�X^Hs�}�ѯ K#*�&������a�����K�͛����Bb��??�~���	x��,����i�[�2nh�*47oq�,`e�� Cb���>MV�#`�(��:$��%ўV)���{%E7g���Sϝ.E�U2z��ާ;�7���-m״�]�*-!�2��H��6è&#=,�� e�8m@Y6��ϧm5+��ß�j�~W�0NHn���u��4�~�Eg큱���r@j�.�W*&e�Fbx�yy���H,"��VJ;1��>;�0<}���qވ'Ϟ�sJ`����b_��B�w��$�^c�$�mc����O����x���n� ��>y)!,�a��-}�-�w��������4����#��=Gf�>_��e��Ȼ���o~�'�<J|�EO��'�f#��!��#Q��˺7+����	�kTޠ�i�Nd�/��N���zH���ȹU�c�W�`)�4|�e��0�9i՘�v��i��`4��V�i�Ϫ(��5,[�=��ePY���&i낹=�W�X�X�lz7��u艆*wO�4�?.;���,8��k��Χ�J~�����}o�$m���
��gz���2is��� K��j�m��q�D����{��j�h_�L3D��
dϮ��颴>'�@Z��d���ZO����KQ�0oH�)���p��^"l�r;5Uc���v����,j��
Vф%��A�y���+��MK��ל)���7a	#�1έ�<Y"Y��k�:[�O��N����ơ��#�Wme�G�5ȂJ�_�J�x�A��x���q�5��%%��a�}�xf2~�M�=�i��3c���p*`��ɞ���{����N�6F���,`Y�0X�O��2A�I/��{5�l+�����qm����x�ָ���C�e�E�1��ڤE��=�$D�[{���M��?"�U#�ʕF��͙E%�kW.<����t��n~:�)��g�q��S:��j:��s�#roI�L���T�Xq�L�Y��J�p�%��5����e���I� d�O2����-���<��Spp��|��j��U��n�tv((>76VCt�!?�p�G_p��~���������7l�Us�n��ɑwn"�N]�4ܕ��5�@�/,;D�����n�AĔ����,�A�\0�<���K����<ٵ{����k��%��\��|��k�7FA��9���m��V�]h�U2U�	ivB
���դ&�a�g4]Z, 3<`�~"nek��L#Y��Mk�Nج&�kI�5�҃����Y����0e Va^��cQ���f˾C����/�E�*��T��TNVh Xg�����)��~��;N	�_����>�u�l���nH�/�րWH r��^i��|X��l)u�3
]�b��g!�� ����&�}Ar�.��0��#������%KI +�Ԫ$RN-Ԁn���2�{*�ԡ3��7`0)�����V�LG�Yuz��[[tc��B/��/5����L՗)�4�^S�{վc�2u�i�4�#��﷒�i/�r�bKhRB��
Zcu������^e7p�Ҋr혽��!	�:H�E�/��y��t�$��"����͜���g���M���%�;۶���wO�۲��4�+�r��X1���HH5��	1"@w2��p$���j궧m��t�>�'���`��ne�vv�*g]�U�$ÝJ�-�~
�`�\a��*�p�kY���� �ʒ���*��4�g��-�1�Dg�
��$p�h1a�L1�����L$ӓ����	ђP��o <Y���QKMX'"�ֆ�>1�(]�Bm�ϭ��}���"��64J_$�R��X��yi^��zw�L]~�����p��~-�>��@�/���u��>��6�Bw[�Bt�DbQ���#3���0<)f2 ��� ׀��6�������62+�M��.lQ�Qe3!*�	�i�&Vx}�fz�f�+*���kݠ�z�lh��J$T:�	�d�.k�J��47��x!��P�����z���S�3ߣ��p)�ՠ��ā(��X���,��!�xx�˲� ���}]H��7XG�̎B'�k��@VHB��Ƥ�x��۠&�����=;d⋝-rڈ��.�<����h�Z`}���Яx`ݧ;����x�~q���@W���Xփ��eeJ,XV�� �ƢФ��q�ƙ��v-��oC��~&C$�Q��OAa��P�6��_:V-���o�������+K�D᮳ѨML�t�Ԓ"H��\,6��g��s�t�)ڗs_���e���f:�D�Q����ϣ�X
��\��R�R�Z1���&�ó�d6�D�|�;��k&�13\����;bT����ǵ���ƖV��̂��I��pk�LY��������ןo����*ܵ+x�������g���U��،)x��q��m�<1'_����i���S��:atZ���ܖޘes��m��Ӣ�t$�������1�)�k�>y�#�P����b�dI,�%&n�CK��G�p$&޼<inm� sj"�r9���C�JJ��p��2��)��d���,�k�C���P�#�>���ԑ/wHrr$���hK�t)�a�&�~���o<V��3��^ ���y�eb�Wg�H��wMKi��ܭ&�-��i�P��.��]����%��TZ�:���2-���rr� +��,G>8�a��u��Ư֖-[�?��ɵ�l�������I��hRɜ���qhѯ +3�jI$X�vL��{2O���I����5MX����5����$�ڌ� �X.��GR��A���%��D!J͘�Ȗ�
�����/!�W������8���3P)�^gwODv���6��4
�	#�nI&�O$eP�H�%���JT4���a`���A\�tXR�"$r�OG���1���+PH�����',�ή^����D U:���S`MQ����C{J`m�\���C���'_��.��� �C�'Ң��?Q`Y^��dbAK%3N�?��'�ȓ��+�9I�Y�8��j�+K����~=�
��]"�.�R���������e�=~��s��g�a�H�IQ]Ą� QQ0�낺���	E$�$�$�d�ɝs�ﻷ���u���w���������ߺ�}o8�������c�	QL|�I4),��bç_���O��h2��:�AD�[��H��Bvnܞ*,]�7���G��[`���Xthz�`�N��)��ǥ�ݫ{�P0�9s�b��E(��Ar�ֲ�+�^�O54&�#KϞj�G=���Z���z������� U�	2N����$yc���*���7�����<!d�@l3	vV���o_ѩ��\{����ӫON��yב+CH��hcjmͰ�^��<�(�6�>_Ȱ.v��ըg��83��=���2�Vc�B~J�)��Ch�9��C�D�^�s\F��C�FEUH�2�*�'�0� ��D��5�o�k�}̞YT�=�\٥��-F�BA�0��	oL~�7l���`�=�D�Y��� �6*���<���3��$2� )����X�j#ܢ1Q/��ON�H���h�|Qsm��\�c��"r�����{��p�IG-���ӿs�C���*��3}jɖ��FE���������f��%h� ����
�<�w���U�V�^y��[~:�;�8a$p>�ՙ�eX<
㮷�P�"������x��x��d�9�1BT���
�-��Uaܽc��RU�>-5Sߝ�E�ײ��X����wy)�l	X�t=^��	,v:������hP���;��i���aA}���N4�� U<��k(��@�	��B�Z�TMlW	R�S��c���	|��gpU�����3�7�d#�>��1	507e�*>�c,MF��v5��sqY�;$'����j�c��9�A����p�x���;yK�!y/�K�Bj��L
B(�`U)Z7�z�Gۂ'۰��r���G�
�-N6,��#+SqMy4K�PP� ��Vu���_{�_W�k^S3&�P����2M�PvE,z1V"}�P����V,GϞ�p��	�yɉ�}x�ŧѨ~>�o�Z������Gs��~���ؾ5�+��{�x,lVļ������<��8ӿ^��KV��vI�KeX��LF��J4̕s����^��#G@����o���D�9}8ڋ���:��i�l����P����<�Z�P���-�4d�h"�7.�0�F�Ԡ����Ad�cY�����l�9�G�:�]4�RE�=h���{���Gm�Z��T�暇B�t5�'�"N)&�����f��e��x�8�y�o<�ʰT�95[�����ʨ���F��u�9_��W�Fzɦ�´��o��O�9u���5W�����0��/�C4�e$۝�f�z���[�)�p�BL���ᵧ�G�zu�xÏ���{\���<.��,�;HP3��(ч�pUc�Ax�u8r�8y�E�ui���N��$TAg*�}�Vu�G�iQ��h���:���٪A���Ω��;���Y�f)��!꣪�̏7,_U)Zf~ңu��w�|m��BEQ�>�F�۲��5~�Ά�:D��S��%:d0Ԃ �a]�c�-�U��j�Qw�Y�څ<҅ja�\'��Փ,�	h�B'�����������o糸�����3Ͽ�-�6�c�x��G�ŧ_p]�ƿ���EK1i�L�@���	!����a�w�vZ�4&>}
��0�K_GT���8�H��f}zQ�����������k�����W_źv �KQF����    IDATՄ�T?lf��:�:[�շظ�١�4??F=�Et���sZU4W�d&TbR�}��A-�Gԉ2�k�c��hQ/�����~[ߓ4,��+���m��CB�f'�>�ǪaX��C�P2;�ڐva�4/�U�k�O ^@����6�u~}K��,��Ei�� (�AgD$�!z�a)�}�\��W���u���Oᇭ[��s��'e��}}z�F�˻b��e���y��X��;�b
>��s�C�A|a:���x���C���8t�$F��Y��	���=K��F�(/+�!���$���T�Lf�[��'Of:� �����C��/D�]��T�mmM�i3]4��5���gA�:W��}�꤀j}����U�$���2� �U=
��
4-H���%9�G����E�A#go�s�ƚ��1�H���E�$��!�XZ���Z'5���R͝C?��bGa͸�|oV�ވ#+��I"!�v�uc�����˱z�
|��G�5k����^{��;c�܇[n���^�EKW��O���[�/?~���l��eqF� (G�Rn�����D��9X�j5�9�=���6n������b������Æ�ߘ�ь���/��q��bFX21t�׆uT��v5�Vi+�j�ż��<��f��3�MTǇZ���K|쩅g����y5��и un�����r�ы�ͣfm�sb�fXDѣ}�p ��<O�jm�Xq�b�o#�ՑX�Z������_�����I��ڳb�M��E�0�B3�N\֩֬Z�������G���7.�r3��� ̜�B��z��pʇ�Y���G��[�8}ʋ�ǍG�(#93�r
�����O� *x���X��{�s�w��QF��3g|ƒn陙x���P�^!v�܇_x�h�^&�F��h�s�����4��R)�}U'L�f����l�H����PX�V�Yk�y����:X}�(tXP4��<�k�����a��d۞�AJ��Q��D�Hzq�"�T��Vê�>qê����@|-�\�����IM��y�۳%�
��s�c��Zt�Jp�mp��c�w�Ƥ)6l������&��u�ݸ���~��aɒux���as�ѢI�s7�~ر�?�.��sr1a�X�$�]���Ͻ�J���Y��B\���{-[^������)3P^FR*NDd"qSX��$���~g͖���5��?5����|ì�k�Z�R��\��Z><�@�G��V�UF�����Q~�M2��Mú�摳��>1H3,bi�,��#HL ~��ڰ4���}B�/�ݜcH5���y`@>�kh�h�?�����,��g(�
�`��#��ҮX�tfL��dko�5��	n�#G�$x���/�
�Vm¤�>eQ$�����������7�#(��W%o�9�w�/�A8l0艷ˏҒ����[q��Ws���K܀&�D��1b�z˶�GTTg�T��8y�֭��qd��c�g�P|Zs�.T�M�2�f$�F�ϲI�U�Fo.��&�"t�p�Ia��N-�'�����q��d���{,�|���U`�,�jYd�܆P�"ϯO�����Y�*��@�kT��j���;X38�Mk'�2�Q$�7���zt��u0u�t�%x��Ǒ_��l݆G}�y��9W������3f!���"E`��ѭu+���	��4`5�`�˕�wߟ���dKÙ
{�$R�Љ,%�8�aCn���f5�UU���FC��ą�������5�~�Y��i�i5HմME���N}ikU3#��5�Fj�x�<N3Y�����a�1IϞ8�|i2r:�B�z�s.m�{������<j�����)N�-NޡQR�������7���� �Ќ����1G���\j����d�4��{�x��`��vLL�T�6�L-�CIƑ��D�$;?|�C���H"=����)��F��Y�c�z�$I��
0��0a�[a4I8t�&<�d�&�*NI2�:b�t(-9�A�Ŭb��@|a?D���K&TT�`�%p׹ڀ�HS�G��8�M�R��jPdX57�;�gi�I������g�P����={,z�(p���l@�S��u�to�wϨ�#x�w��i��R�0Y���b)�$s%�}i&���������"�8�U]ܣ�T��u�zRs�i�,��V@�>���B��~$'������ݖ���D�"D(�0kQ��z�p�k��t ����hު�8o{W]�7��:��z.,[�
�*;l�ې����?�易����e�#BJ�3g� �a!�H�_]���٣�1}<2�v+TOǸWz��&٣1�J�i�^<c���0�[��-�)nZ�L���dXv�6���b4)L]|Y��1���p��G�5�FM�~�h�'B4Fv&!�f���B��>Brkf 8+񦓁ir�n��)��CO�ǫ����xq�j�	TK�J�^.I�;�ܤ%.S��E&�|��N塢r�ژ�vq�r�"�=��u6z(DzACzm4� m��z5��|�jv��&)��Ç�{�.#��㯰f�F�z�jO@�����dRZB�(���G�?�6('uL�:�Ƅ�;(NN�N���q���L�7�	����gg�)nl�HS��D�$���h�N� �*{��h�x�G�gCx�� ���@d3R����u�r��z��u]԰��e���sE-�vm�z;q�A�U��Q�dڌT����@#rL졊&i�~�K'#V8=u͉Α;LHUM����|�Y��s��m�H��z֨L�<�'�8[�{�ύ?8nsq
�8��^��;T�"�0%��j�������qX��fOGqq��D.��h@��d��ړR�rI��נ�TQ��Pѫ����ik��w�(��7��ݨ�Q�<�91!��y��Fb��Ľ]*��b�(b�Q�����r��U�!ݖX�	�`��������F=�lo��N�]��\��K[f�?��_~Ӱv�?5��B49������c2��3�bAb�[��E��\��*ɩ�"�dZPr�js����2��By�h�:��T�C�ݣy,u)���C9�Ҩ$5ާ85��t�R�q- �jG��i�!1��I>(ۣr����)�u�fi�>F���Ph�#���0@ΑB���0���h#�r�ȗբ����EG��H�c5�-��S����&U�'�z���67��h{i�d��h�A����3�x0�?������ne��H��eg�F�
I5�0۱�k��Q���a��i�;���U��YX���7�t�S�EerYIG���/j���m���S.�;�[�1tjn2F]�/�[��'����� �q�Qi��5���g���qAп���R5.��k���>Ӿ�qd,�����o�8����?�`BD��F;����?0��{��Xc���h<��/ט��%ь�����pTЬ��T�{,��	b�&�gj5��Kl��KN�3��-q�u��"�3҂�?1A�t�t���t�J��q���<�oV���&n�sr�N��)L"K��v�o��j�����d�T�3�-�����z>�I���yD3�t�t�G����C��sy�����rk�=�G�pY�V<�bO'��q/Y\_C+��|���q$��Vy��sK�|��d�s��2�c��d�gbģc�tq	�f3��Dĸ�����:'��٩�U�ִ<Z�����̨V��q�%��W�^�8^J��W�zT�"<��Q���}K�kW����u�����t4������Ln�'!!�M��JI�$�b�V��3�ׅ�Y	kz�ͻ{��~��Q����/o�}���`�"�Y��ZH��@a
`�Y S��S�b �>A�H:N�S�/A�ťe�<���F����
�h�,�M(W���q�jNE�Lg(]�R\�vE��yL.���/d
qU��:�>�JM]&�T�oqo��,�>�s�Eh��zl��k���šH"��\"a��|lP4�I� �si�g|��X>}y���;4RY�ԊO)]ذ���=:�]�G7�LF�#��%�,+iB�L0 ���R�*Ka6X&%%��as�PU^���r�����?�jbF{2�� �P�����j�
�ܨ����{�����5��E��-c����ѧ)+�Y�RR1��M(�j��ݮp�!���ѪY�i������
8z�$��*ƾ�q�LA�#z6.��U��{g���EUmD��w�ʒ�U�c5X�9N�H�O�V3,���g<�a�'��K�
Yg��j�*�6I�Ni�X3B�r��,�²�V���#B�]��T3V�>�����FI#�ijΜ	�@�C�ܦ�r�o�qiD�"�n�!��>�
�J�y�}���__�lՂ5�	�I���)��=V�w��g_���u[���EgaE6�����Ib��Մ@Ud'n��,w����a]{뽏o���UA=�MŔ�#$XLH�ZQVr��-�6D�+z��3�ߞ�JΠhGӱF��D���(:S������t����l�#JZ:q��|��E;��G�<q�k���y��ϲƨG�JT[���TM�ҦU�� 虒����\U���>���璸�v�|����
1�>���HHt0[���CD������R|��\�j�gU=�rXT3d�c��L�9�y㩅�p�ؤUyzv��%X�#^�8�:��u���|RL�/���O^|QL8�Sŕ�;)f~<�����#YH4¨��nF��A�l��6�6nؠ�5���{x������I�J$]F�pv�3쇁��a?:vj�NZ!#с����(I�D��Lx�F+��cb�{�Ɗ�T7�^�4�&~�Bd,��ś��s�:�aϥ҄G�c��@�2��1�`�jZ!�~�V�U�:��"��v��;D��2gG�F�CP9��LbB�J\��8�=^7¾ w �Di����1���l��GHh�x�jIaUo�#����j�<��'��Z2!-nu �jM��:H�
�S�N}]j'I� #�	1�G٩C�Lq��Qw�u˦<��{8{���c�����M�r�k�vg�	),������Ù_���2�d�q�b1��v�I� ���;:\�2��Q�~��a�k��������� �P4����dU��+ѼI#\է'�S���}��|\��̉�1U(���4�J!$�5 ��,�q���֮�7 Ö��L\9�j�V��k�{��[�GI�H+������q�U=��!DU�s�e�F5�*�Tω�p'�$����T�����L�iQѤ4�04�K�K*>�=^n�P���/�\�3���)Qh����7%4$CMt
��C�\�cE��G?m F����\	'�(����=�A� 3�	�E����KK�߮탮Z!��/*���F��DRu<DB���T�a�Za�%����i3�c��q��9�#��LBr���"�I5���(e�c������u��MX�a�� �,�F�:!�L�\�$�����Cǖ<ut���h�T$uU)�<)Hq��`F0�,V̛� ���lH��Fñ"7�S$ep�U����=PF�j�5hذh��3$���q�
8�|i��IK�֐��,�6��&#㽩=���3�fG�D���֠iLWU��\���ɱd�jA̝�i�p��3�M�P,�z*b�a��@21���F6h��ӈ?m�h��p�ϱU^f2��E�W��A7��~�`b8y�0K�)�)at�*��_��<ʒ��88?�1J*���;3��W�aLȄޜ���f�R̋���NM�F<q�ȵ7��_�a�$�L�_f��F$���(����F��+a��*�D�-��(P��5���1G���GPeׂ�R|39���X���tTЏDs���΍�	���K�*�MBĹ@���b�!�g	��ZH��b��P��鸩�'��s�0�W�&.+YHj�1�Ve��ܮ�,��f��~YYq�y�����u�#ƍ���yhD>�-�(S7���5�-|$��Ԧ�"�*\�G$�p\�Qf�Y�UD�hR��GǏe����^R�5uH,���;"S�p�j����lg��e�v��_���n$����Ê�r�9IҁvG==a̪�֭#��|�Ήި���V��,+B�E�>=��k���y��0Y��S�����ؼ���0���Ga���.^�U��dNDbJ2׍����Q���PO��Dur�b!fm����e�$�ĊM�ARU�)��D��j1��S�<�Fߙb:F�BFi�HǕ����t���ɃQ�^QZ��Űbš�P��0��P����E�G ��oa2�����1�A�LL8�s��悞����AR��ȣ��"a��S�N��I#b�*���Co���x-JNU�2�bvZ���W���B2+��jم��t$�6�/,��W�����ӓHC:o*��N�o�:��F.��a����k�M"�2X�p� Ѭ^؋T�	�ꅖ���+�b(Ug�x�2 �~��Q�����-I��;��>��箄7�g�"���Ԟ2EMo�]=	K��|�z\U��el�Dx=�jc���X�|��C��> �j�v
�{�|J4���*�Q�:B԰�!R��P�0%�u���` F�	N�X%g��n �a�:�d�%�PD=g� %Tz?	�i^�2M�(1�m&n�W�� ��H���;k�,<	D��ҦixDdJ	�E� #������x��	�ت)�N��plH�j��6�Y�T��gG��$}Gɒ�tVi���:����gp�'&&72u��7N���	c�u��+/C�=q��[^�:�ɞ��4'��M"n��Z4(́�_�JW�Q���3��{n���Ѩ:�M�;RMp�ʏwg-��7�2�`�'���0&G2q]>�S��BA��r�'h�Y�v���UI�N"c5xG�R�[�^����d�!�ޅܼl�����py�v�'��`&6��i~,�L�d�T�.-9wU�V3{j�P�6ǁ�G�#Ā��#��5y �Z�����A�|npWU�A���M�T��UE=2s���_���jJ�R"$%J�1�X�	&x+� E�x��'Q'=	����@8&3�ٸX3Ѡ�	,�b�ě��()��H̓N?���z����x�p�Fbz!#9�'>#A:ܱa�O?8�Z�W�5����[���]!,	IHJ�#����"�1�[��B��R��T���|ψ�����,��H*�_E�n �,�<|�3�,��#EH��KLE��C/�* �l2B O�.C8���d@���e��
/�È����ƉSE��{b
�4�0(��8����ѐ!�IN
sY(�J?<�E刉f�@�3AOr������I��<aʊO� ���ec���DVN.lv'��ڋk��ޒ�Ĕt�.�e
4�dHN�� %���4,-�7E�u��?����§�}���Cf݆�&����pa��dr$�}�D�����G�h^�X
<�
�j☗�,c"��j�P���('K��D�DoDR�J:�9��v�:L|{~9^gz��Qu?ө?ܶq�O�?��5��g��]��`�`4#%%r�c4�T����c��(>����53�Y|����7��c�Ͱ�s9�X8�|
�K]!���b�>\���\�ɣc��H�g#��v������Q7lF	�pK���W�SP�j_�:�Jo�%f{
'|�s;�Q	�]vR���nB"M������Q�^#��
���%U��d�Nx~j�F��`�Yp��!�$d���l���QP'��\�������I,\�����L�J
�:d�X����UE^��C����l6r-�k׮h׺	��8����v�59�����1q���ce�8�H0+�W� ?^|�d�$p�E��R_���e*��y+�U��F)�0BO�7��F0�AVN6M���o�?�J��&���H���O�n�8㞇���Q8l�s��_�����`tezF¾
؄(�R}/��/���c\"Uu�7�"�|�\z��*(�#�D�5�!��$%:�������R<A    IDAT
=�BJf$��f����%�	6f����:��٠0���?��0rs� � Yٹ8S��O����v��~�-i�*�r���$#%��C��	(r��N�ׇ=9?.âU�5$��3K���y�JQy��fn�ڬ:$%Y`�0Y-(���сw��=G���9S�jM�\�6J���I��"a1*�d����V���r�\}��نWޞ�򀄄�l��� ���� Rd%��A�_�ƍB�&��*;S]� .Q��U����,г� *��F��C�%zB�Y�pe��%�L�wP�5���)!�I5i_?k�#�Ͽh�>b��]�~���;Z��!)H3#?##�ݎʊ�\���j����Ү��NP��eb�H��­;�����!!-�E�C�wQǡ��Q��u���j�aB�{ˑd3!++C����>��[ɩY8Y�Ƣ��鑘����J�.��?C�`�B��233�Ч�d�����ȭ� �h����PqL�48�x��L&��:�:r DY@�F�eُ�yYHJR+�z�$������'q����IO\�2�VLb%�w�^v
rR�8q�g���s6lؐ�>��^�:[c��-X�y/��8C!�_�H!��2C��$a7\e�q��Wrq4	����xI�;���W)�IT�N�o��
9J�u�V���31���
�%�YP"d%I�;6�|��	�f��a=����6�#��-:�u1ȾJ�:ad�m@?��Aee%S&Ү��8U�)m7�-��AI(ã���JF3_�h�Z�]�	z[
0G�>(WU�䠛�ղ��@;0J
��w���
:r_ϙ�*o y����mc����������y�P���1���"���UW]�;߂��a����K��_u����}�qA�h��?�?�����Oe1�~:�o�˻w��ӧ�u�.Ȃ	!�PT�ŁC�t��Ʌ�Mz��:����QA�lX���O�=z4�6m�I_Ů=�0l�#�s�^~k&�IY��j�K�d�Y/�NF�f��(�Kø�#���|�Y���&q�2�^ D�|н�z kk� � G����f�
L��k>U���6Q� �)��� 㑧��Ӌ��><o��WB���d�`ѫc�&!��9)�]o΄<�~���%h�B�vS�
zӋ�5f��]�G^��;�3f}�-~�w
	iy0Z�R�F�(�W�~3"!�u�:���n�E
T�jѡ}�1���_�~zN>\A�T�a�xL�c��:L�a^*Ĩ{vm���F���x��'PTT��?|�ehݥn>
���;��3�~8�)�%����c���>ΨdQL�$���n�~���8S�39�v8	_X���`Qsj�����Cߞ�Ь�.6�]�#�ra�ر�M?���$|�x1F?�����ɟ�`K�՞�8~���p4 �B�݀�4d_�������ť���"8��4�P"��N��Foҳ��(3��j�#95�Δ���_a���p�t�L�83����R�v��|���_\԰FNxK6���B�Hc�`�$!�b��ꇙ�m�W���@�����jY�U�FR��p���"#�v�т��W�e�p�$��0��%��h����$�81Be�QV�9X������C�+{bǎx�ſC��H�)�;$�ة
�b:��)5��	�J*�J��c8~�g8�\wM�9
k׮�˯��͌�ݻB�9�e�/ض�0̖,$&��2���pX$[MjF�WСm3r;N�8��k6@��y؉�ŕ�}�9��Q��+q�W��]�i6���-���6m����y���p�T���gt�s=���Ĵ�!(��Q�yB9��¦�u���MK�?��������.E����/).���l1������$���7�@DeyNIM�39GN1�a��p��U:%F�*�/�H�	��5H����5���x��a�	�si�>B4��$�Qu��]۴宺��F(H]�ۡ�w�I�X��K��ԴL��{��O?a����{��-&R�⪼�"�nG�Q M���N��I6�0��Z^�����Ո]�va��]�%%Þ�ű�ƭ�Q���	V������TA�S��d��$9���UhѢ��ك�+W !%��4��k�G�9	΄<Κ(�LN������t4�f�-ѭs�)��c�����		�}�$~>v���ZK^���)���?�[�KЦI=���U������	�
��6@F���h�2,Z�:[*�Ss�r�<��r��B�!�$IV=���A	y���@�^]���l��	wP(Q� f�2
���SE����ث�J�/\��뷡�< oH�+���L�5!�Y�(��tꎷ������\<��Ћ�.�~bPtBoq��@"��(���	���@,�E�f�Ы{74lX�����! �@ U�uF�mNx�!�U�����X����V   {/8q)Pk��gt����>�L������d7"-��G� �����$H�#)Yy(�����*+�@ J3V����JuZ�.;���-��CVj"l&��*/���FE�;����;�x�Fk�K�Ф
��h�Y'���hBZ�VиQ]�%'0���LBq��vGq����T�����Lb��c����|#n��Z��n �U!�a�z��-��}�p�#/�De	i��b�?LMl"{-�!1(!$��H�造���NZ6o��W�D���z#�6�A�,�b��`5rkl��X�h%v�=��X���z�	)��=B~d%����>���w|sQ�5��W��d�?�$ `���.i0[u�
�b��Rg�����(�ָa�l�u�Nt
��O�����������q9V��
���"fJDDTU%4Qp�{���c�[��S\�uq�#�nF����˄�b����dxɁ�Ǳ}�Wx����(�ZN����<�NO@��u��N%�,����4
���w[vdOC�hM+����9I^:�-�^4���Fu�Ѵq=���q~9r{Ɔ-{�[��Ѧvu
,:�p9�N��K�gc��p��}9x��+J^hl��vb��X�~��4�2U�X�^���zO)8���
�@�+ѩ�x#*� tRi�ԯW��M#� �Ij��LI	>������YM����Q�Ęm`"���mϖ^�&����O��	w}{�둉,�~�7fC�5���Ov������N��Q�;��U䁤v��7�8��*���GY��.?\�²�t�z�4��Һq96���+@h�U3y˰O/ZvV:Ru:#A��?��r<p��I��a�MN�vƃqr�P�C�cO+�aX�
�0h�u�ݧ��_�E�Vpi��I����L�M�IaB8�նU�� "�"�:�����:�LN1屓E8r���}��@����D���8`Arf+O"�;���$t��
�4k̍���r��]X�~~�w&g.�2		�$�T���h��Hr�����H'�� բ=K��&�)��6Mިx6Z'���!"��p�`��J$�1��39q�Y��W�� �~�mô{���E�
~u�w+7�����#i�K�F�B�êl��`�!&:�Fn���Wm��hr:&��s��� #bn5r��+�<�W��O�poP7�Ԁ6Ү�	{y*���%BC���e� *� ���G��3"����O��#��9�bn�iw	:u�5k�a��_`����#�`Ic�*58���2��l3Tu�zOs�E S�%��Ne��,�@�,Y!��@�3{,�w��0�d�9M�C%pU�BEe1��:xU`3Z�� ��9a��'�Өs�܅��Åd>�8���Q<��Ϭ�a�@OO��f4�rOPO��(�����E��pb���$�cb��d��b1�f�	T�0�z�]�̻u���C�hͶwB�����T3V�gR
��,@��.�4�N�%�l���0M�Ќ��}��Kd^��^\҃*�ŇR�A	*_XzD���!�<4aR����i!U��{a��z�$廉/y\�(i�6��(�q���P%BAC�	0(Hf̉��6�����)k"z$��"��#���g�:�++�r��T��6��3'����&�Tx2t�ЩL`ћ!MT���| ���<��:Xf�	�Eup�ɣS/�	�5�cI<�x��h�/��h܀�=�>�ť`�R���O��	�D	ڣC����NFy/!G�ؖN$���YB�[��L뾶��C{�5�1����������)z>�
K�MVM���,ԉ[�3c��$��
����0��'��Qˆ!��60�����9��xk�周�-J<K�O$������A�f`z8$��_T���"�0Z<�Le��8F�[#��"�SFk��C$J�t6���P�*qB�JP��i�H�t,f�D���Mӱ����EYx�4ED=P��Ǿ�-�"�H��Dj!�>Ӄ�"1#\E�43`��	����3�&�5�������b�Q������u�֠a�֐��u>!	'�ܧB|��9z��f��\�&�3�D~�eoˆ�?>b����}OL�n����?�?�$�*ɟ�aiHKY �&u*�0h��Ӡ�<�̼�q�L'�G"�IZ�-��ş��S�"AK��v�vO:#Y��P����~������HIA'�`�� �iV�NG��H��^e����F��G6f�0�t��"&ze$j�H1&�=���#����h�ӆ�������@
�	9>C�)a�������c��3�P����qFCP�G�1��R4E{�n��o~�ٱ!1��g�3���V�ɘ��RgV[PL�MY�H=E�z�z�`�2,���O����w\|`����y��͋]A���@���ƌ�x���S�_�?�6�Ju��UQb��8�${ �k��K�,��Ƹ��Lj���u��N��O���6i�[�AP/��$D���-�{��3��P$��~6l�р�h�����Ltp� D%����9Se�%�D��9�T	HH-�Ř4&��F����JTF����I�H0�TL�	�Bs���� F�T�R=���x°3<L3��k5��5rZ{un@�gMF��P�֎��,�!9�1�J�'��}D
BjeF���0�߷��8�1C.��E�I��.Z���J:�@p��C��.�X$*�� yyF]��T�E'�ׄADAT�T跨<�J,*+1��Y�`M=M�����A�GeY6���&BRhA(�Tb�Ng0�F�^��ubEE�>��V�]4��X,a�a4&GBaQ�$I�ɂ��b&�����c1�� %3t�Q����7%��AD(�aO�~?�S�F�G��:�Eqa���*m�,��'�;�-�n��R�H`o�2Q�lzE�	��yAc����QAb�qj.G�/����j��X^�*���zc4�rL2�c�)��7(@�Eb��~^L��L�h\�%�?Z&�C�.Y�ߟy���BaG,�Ag�E�J�^uz�$Q��כ$�"I�l��%�)���Nug>ӣG��節~��'���G���,�1��3�"�bQ!�2 ����3�9��bL�	Q�u~uQA�����X�Vd��bQY�
Q�C� �1A�f�W2(�()6�5d1����g٘��BP���)*ʱ�����`0���R��M�:2W�H�MAg�%%,����P Ag0�}��$%��z��(>Q\�h��u�3�z�y]Q�)QY�ƢE���2:�_EwL�mr4�0�L�٤���c0$�&��>�N*e�hBVbaY�I:IW�Κ*a����ɒ^�b2�����p(����Ű[����/��gE�z�6���)zJI&�	�DA�J�HX�E���ڊa�3@J��3
 "IBD
��$(���(��H�bĒzoN���G�Rϧ�����k3?*���)���5D�k���_oC�#���y		�m۞��7Z�l���{��Qg�L��Q�$I���XZ�%2p������	e��4�� 
�2�t���fumע��w~�?����a͙3'm��M�VUU���c�뮻��Ts���]�j�i���,�p���L[��}�?���=���̸<��wj��?b�t�w�M�����6m��f�=ѨQ�j��?����|�_ް��ꫦ�/������G��[n�����.�o��߼e�Ċ�Ҏ�ٹs_z�񱵽�v�ԩ�y}��~�Q�F4Q�WQQ�勯��T�c�ԫ[�缼��[�l��V7��/���s�,��h��f��Uxn���X=��{��������/���������S�_+��xM�<�%����+�ӢE�#��ŏ?���t��f��K�����yw4m�|^m��g^��7���5�����P$���*t�m��p�����"�wqg��沵k�|u����º?�;r�e�;��kϞ=���V����sX�歫�~�8�2��9KEQlոqc���[�4i>����?���Z���/?_��nw�����4xȰjP��]����r՚/�%�+�����o��iӦ���~���b뼹_����.��ux�6������)}�eKcr�y��]�9y�6o�zMm��g^��7�-��՝�٧K}O�7�����!����������/�Z�fŬʲ��F�o|�-W���hϞ=��W/�B:w�4�M�N�6�~�)}횕�B�`�ƍ���f_޺i뽿���'\��7����gM�5kYyiY�`8��߿�ȡC��:���z/^��S'N85j�e�]w�hѢ��j�"�5�7}~_�n]�oӦÂZ�  ���+Wʈ5���;^�a�^��49X�������k��ԩS�.s��-|>��O�>�F��Am��O?�l���E�N�7n�y��^�977P��PF�`��K�~��]��նm�Z�{L]�d�ZY��d�mT�A�K.��Zd����ϸ�/oX�6t|8���`�mUUU��=�7�]�i3>�x�Y��Ŗ&M�����1��ׯ��}�c}�ݼU>��n�]���<�K�.�^�z�Y9'�����������w����'��*�v*++w���Ə��a����^˖��_RRbjԨ��{G��ִiS*Q�מ�=��6n��=�;u��S�Nsj�v�t߾}�KV��"�bAZF��zt�?ê�*�/����w�Z�������]�v�����Q��N��р�˗QQ^�kР������x�C�9W�^�����w��axǎ]j��ٳ'c��U?������z�Q���Z�������}��#�x��K++˕nݺMx���_��Mߛ9��U�W}�r����
��wϘ.��E��jՊ�>�7�]��#:w��am��Ν;�V�Z�U�I���ig�7jԥm�f�H��ߟq�_>ƢE7n��Ғ�>�5�~�e�x�Z��~x���+g�=�7���ޱ�v�#�U��}��5�}nO�v�;�ձK��k�`ɰ��\�E������Ӎ4�ڼy�jɶ���ϸ��°{p��GO�����C�=&����j����}���+V~J|�
�����u�ܹ�Y!��������mݮ�m]�\�um����+7�t�:y�9��/�ڢE����ϟy��a=��O�;uquv����Gz���.���s�u릓�����;ꮻڵm�V%��ŋ����[�nuS׮]�9�~�m6��S���oJ�:�s�3��׻�u�������	��w��||�T�mD ۪Y��x�'k��'�=l����'���ܼ�cGk�G
�G�1�\�r����n۶퍝:uZ^��yϞ��lL��


��6)��ma�����3���0��{������qI�K�zṧ��2y���o|��v�n^����tN�8a^�x��ϗۺu끗^zi�{��7��X�t���V7�0C�����k�����+��7^�����H̱~��������v�^�<u�7N�UT�NN��Kҽ  8IDAT��Nhݱc}��/2�E�m�z�mڴ��{���c��6��oϚ�`�K��^VA޺����������/���0�7'���}?=������5���^����5iʴ'�l\����rr�~=vL�V�Zŕ�~��6�aÆ=qú�{��3���+�nݚ�r�7k	��9vԹ����FZ��s����W�;Ӧ?�y���B� ck^z����j�H��|[6>\Qt�ٙG�=<�M禝+j{��/^L�U�m۶Cz��1���شsSΪ9sW:��y[6l�������o�~�G��[�����ᰡI�&�_yib������za�捏W�BVV��Qc�w�СCym�C���˗��}��Cz��Uk��j�֔����lw�L��XֶC��H�����y��ǚ����-\����h�ԤI���=�z��.��S^{c��M�*N������n޶�m�31B&,X�`�����ԩ�m={��#u,��Y��ٝ�dfdu�]����������k�֭�]%{=Ur����	������<�w#.i�jә��,V1Z�f��p�a�����kU*X�jUBeee����ddd<ݤI�ٵ���\�$�h�w��&Aw&$gLMO)ܙzm�Zf�Y��6�e��:��X3�T��ۂ�`A��Ѣ'6�_2�	��k�r�m���ff���;O�y�x�bhH����8Ä鶤3�I�t��4e࿨��ܹ�:eʔv��q�ѣG���myyy���uu��e��_�|�޽hP��K��5KǄ}�}�H(���d���r
�m�vN�~=������>�/kXO|�~�%�>����zz���tP,:���A�Ɉ��O�%�{��ޣ�%ek.���>�"�����g�DP"
�Q�"��wkX�5�%�����	=o�y��|��7����'lڴ�{$1�"��4�G�AR-k��ǌ�#\�^~9ѷy�åxX*�����F�E=d���/|�ɀ��v?���Ai��/kX7�̼á���� #��Q�Tt�D٤93��J��g�;�M�	�[��1�o�j�j��[,���2���J�V[,�@".TD|142&vK��C��Ϣc��g�[�p���Y�YL���`,#>)�F�\q�s�,Y2P�S\�(f]}�K���M
G���)�I�P��Y I12���a�7�\z��ֿyF����[���-E�ND���P���k��������/���/~�n��j��%�[z��']�ȫ5�ƃ�_}hC���� ���[^�X���f�;�O���~�Гs�/�U�lC�L%z�6���ρ<�5�)��$	�H$"�~���:��=z/\�0uΜ9�?��çE1��ؐ!C�2e��/����#��c�!9�ӿ��f���0�\Y�i�o���6w��D� ���������֔�G������_�c]3��׎���ЧQ�a[�5��_:|��Ϯ߿���;��ֺ�?�x�`m�}��u�����۝��]F��p�����B�{�Q�k��YydG?�A��p~uC�v#4�%
�_|�U+֭��K�M7���'�|������[o�0{����a�k׮����{���y�]��ڻ�Pď�����g�|����u��/N	I[�|�����'�']�3�77}☻gâC&_gCe/^}{��IW��,��6�㩞�N{ж嶂K���qK���K������ue:�-5h����ݜ�����`N��͜�Wo���_^�Օ��������>}����˖-��ѣǯ*�.4^}��Y��YYY����K���G
Wկf�L�5������F�$sd�/�	C�\��?͒Te7��y)ۻ?0�O���J�$��͏���C_����b����@�M���|댶��m��X�׉I	r�)�:?�O%{�����^��,����N}?������q�rw�� fv�hܶ�S=Gr��\2~�}k�`RQ�@��Xi�-z��rڴi}\��I����;���}�_�p����<c�ؽ>N�8o(�h��4��ر��������f&��i�E�r�����9`t���
]���.�Oީ�@FF4�����Z�۷/Oݼ�jz��O�Y[��eu=u�ض�m~9��|�����g�GBh$$_٤M����ʟ5gΜ��Ʈ;y�t�(��U�{���~�7�|�p뭷�������3f��z�5ל��m����=O�����<�DR"#�M/�{}��嗆�C�WZa��*ȭ�2at��Cβ���}���aї�;���=CD�����{���_�#�vM�l��II��h����5H[�/���M����"!p�?����/���-n{���Цi���w˽�\�@v�Х���cwϗ_ƽ��7+6��k��ѷo���⋧Ͽǐ!C��裏&ɲ,���k��/�|全�����S����X�N4����M����uϭÏ�\�/  إ��!���O2����/iXc�zq��%���E(့g�/]��j���v���o��}p�u+�-�	��I���>����nx����_�tߺӻ_/IT995��v��F�R�yۏ�~n����ǖm�4�T� U�DGs��)�<v������7�z+��~r�رcz��9g��%˖-s~��'�͜9���z���뮻��2e�'�V�r��K�N����ϧ���͒ur[�����ܹ��O޹r�,��L��2�L��a�fڣ��d�Zw}��;'<��2��/����X8�y߾}�N�t=����,ʬ�����Əv^�ɽ��)��&������3��<|���32q~�
����A�O�A�Uഏ��[�!j��0�:uڴݻw%��������t��?@�	tp,˟?�����޳gO:�f�����G�'H�r1���t9�?F����9XE�~��󟝅�'��^U̶]��`*��d�`�Ιg_+z��!�=�o��Y�������������':|R����W�d����L�;��r�s�O)o�0|b�� ��
T�q|�ˠ�)����y���Bw]P֑�����[�"s�޽q���?u��������hA\\܂��t�9��ܳj�ė�GR�>�(����t���٘�2�g�$���ĠB��e�W^ɻ����l�Ҷ��ؗ�9������>|�j!�ǿ����Wj�B&U<�d��������������9X~��(��U�S�t���NGm�F9z$�_�x���իf>|��翧��~A__���)SHZ�'5��߃'����w���)/�e�#*+]�O�D�B�]C:a���Q}��фE�0�6�&����h¢}�HFֈ�v�{ �ߧ5��    IEND�B`�PK   ,V�X:�I��  �  /   images/65cd5dc4-66ed-44a6-97e2-8bf96ed14d67.png <@ÿ�PNG

   IHDR   ^   �   [�7@   sRGB ���    IDATx^�g�e�u&��x�=�ܜ+CYI �[���n%$aD,*PH�7zH�����m=$ �$$��L ɖe[�H� +Y�n�'����Z��F��{���FJ�N���s�5�7�9����WA��W���R���JF�o����J�+}�����g�{@�q(kH�����R�c-*�V���c5����ݴ,�R�j[�
T�Ď�$�R�I�"�mY�eY�#۱,�rl��?��X��F�\?���M,XN/��Nl;��45�I-ϲ-�J�_׀R),+�ϳ,�_�"^znj���8�)ˎ�)�4�S(����ہR;�.�ۿ���]pA��z���9������|������/� e!�@h뿇
�,��%���y/ߦl�hi��ߕ��2��_����`��=?c�=�e��Z���"�{^�r���s})�!�3\�>H�$l�[�o|��k.9�1��W��?m6Ñ���c��Q��bAԂRJ�R8r�),�bi�T4`��ϛ�m��s���+w�.�Z��Z|�~��/���GXr!�:,�p�(i�۶J-'M�ġ5�������'&���m˱-([�J�T~�Z�~�)R�XQ��p��f�_}��������o����J��\�F�o��z���MJ��I�D>�#J`;b�D�vl���m#��G����A%
��!J8��0����hle����#��9
i����Ba�u]�\Nq
��`�6���;�2�Q�m8��8��`�{|Ǖkm7�����^x[��Z���D��]G�RA��h!,�AbY�r�x�������?����{3��I�[o��؎��^��G�z��}�0�J-���h���²}�$�e!Q
/(I`N+A A�i�|;�,��s@�W���9��Jm$q+U��B�� ��T���C�E��E�V�-�D	�|ql|�J��	[�ȻlXpr�*I�~,�Je���rE�|�;W±b�.d �v�n%�<a����>l?o[�s�o~�ͷ_�ş���z���W�z.�c�
GT<�����k����	~(V���m(���sM*�s�F�ܸ�p=*I�A8�7�t8�a�%`��:HS޸m�p���t**M��n�q����x�J�������A��%Z
��vi�B�s� T�\�)\�&�`��]G�����o���O�j�ws��3X7؃+>�)5�i�>kc�C�7�^3t�?�O��&�?�w׬�����zugt��;����{P�e{h�cx��-��6h#��!��\�ڪi��j�?W�ޜ;���X.\׆�(4�(�b]�V[�=�w�r|��h�X,��j�������n�P���$
��#P.r�"f�pG�H1ڔ.�GΥEH�&���(@��<�Np],���2�T��T�1�b��n\ú�".��?��hg����#��}ޚ5��?�k��ͅG�k`�O/���]1������	����h�Xv�V�q��v�E�������y2rT" �/�ٗ_Ə{�����c��#
"x|8n�$��wN9'<�-E���v�x����ǟ���$1�q(�fs��c�yG����'�@�݆_��B#w�>�߼vH��{'W��N��N-	0�[�����F�R�\~�H�/��}��G��b�GqE����Uǆ�|�O�f��]�?����?wú?��`ͧ��9e���_ܽ���Ќ����	\��ۨ�>|��8J�}�*��BXq�{���yg��r^�&��B�������$p�<r�p�6Uǎs>�S��npK�IL�����m���w ��z"�+"g�@�B^��#��?�8�~�:4�1
EWb�����~<��s���s�
��Uܤ��6��㻶b�~nCj2ڟm ��/���;�����#�R�]���1\n���X7ZHcL<=5q���|X���g�x˹��q��uD6p�_�Uw}�$�
���}E'Eژ���N�<�4].�A��݋�>�c\��nN	�߁V���8I�5� NZ����>��� ��Cƒy8~���#������Dn�p`�Mtz	�`���3N>�(����r:y|�����@��H�$�&	r̋�El^ۇ�r�Vl�G4�Z6�B'C���*���M��9� �3�L]E�,�P��;n���X?ZN�b5������=|�?t��_qѮ�;�����o<�+��6�|7
������`�P�Y��w�s?�\҂��%�˽�ޣ�����P�=Dn��C�0gT@�B%X�,.��a|�ݧ ���r�2B���'��;���+j�l[B=.��U�PكӞ��~r7~��c�\�CD�,��T>.�~/���kh*a�Ip@w�+�ς.`˚n��Ƕc�H�FU\Mh��R|��/��N~�����"CS�j���1�������\ߟ��?>8v�kG��a[����=�;w�2七�����a\u���Js��|�:gx�����q���� �1ڵ9ٜ�J?���3�����Bۆrr0�NT
�e~#o����������A}	|��^���S����Ad���g#dk�pT���j��s�I�t쑘�8��ׁ�.�kn��z�_�B��/�j̹98q�4�i��O�>GoA�:��w��������7�Ѓ0q`������B�U1X����	l�0�����3�w�=�w����[�{��]���ϻ�����#�*�H\�a�8L$�b\5gq�{~;?���E�/Έ�����֣���ދzd�g$q �w`96� D)�>�8�=�^sJ��Εx���c?����[�0ӎ�H�n�KE�Zȩ:�����lA����Rꑃ+�|y�Y��.��-�&���c���y��O\x�uC�"{���t��<��W;$���$	:�E�v��5�M>������6D�5�����[���d5��+vﾽ;�ZzĻ��1\��{�t�������,�5q¦a���o���Gl���,^zuO�f�<�s$�����f�x9O�ٮ��q�`�s�:�y#�y�x�����L�Ǟ�5r=:���y.���g��D�?�q,6����CWw{�L.����?�+���"LSI��@��)0dѓO��q��;p����X��O<��fjx�_al���ac5�Yk�b�FԚ������Ob���dRa����{��9���O郷��{.��r+]�smg�_?����.��7Vp-	��H=;A�j���w�����Ə�z�߶Sa(�^�&7Cf���giDi��� �4��4>~�i8��S�������v�FԒ<�[D(�~`8h9�/� ��U<��;'��d�~�����/ @��C�q!�h�(�D+Zq���E��u���'��م�/�
�kP�N��>O6]�H&k�S,�H���ܟ�W>�	l\ۍ)`�῟�k�����-��o}�����b��"�����|Q�v���ka��t2�F(Z1ri��wo�������_������$��-�1�l��*�kU��<\/'7�Y	�h��\���x�o�����?Dap�[Z��B�J�l֑�y�#�n�΂�(=�s�98꘣�����C�?	'WAb���Z����y�r�S 
Z��[����	|/����1����p+~��Ax�4�r�خd�\��w+���X�Op���	��ys��c��������6�p�-�^�m�7�<{l����qãϡk�	�3aƙ�!�V1��Q�l�qk�����|U�x�)�ے�����pEc��9��i@{oݲ=]%L�����a��0ӈ�Ps,Vܐg�*�6줅��q9��7I�3=_��Ԝ$BQB"��d��+ƆcNԆ�+�dp������,`lf�R7�a(\W�m)��'Q(�ړ�!��|�|�q 3���c���;:�����7޾�3;���`�^�}�)���C|�;;��
�T�9��L�|+EҮ��E���O�_��.v<M'TXGGї��
`Yd1=�^P���a%�$;!COFvN"Z(��b� ���v$��ȓ��C�a��
�B�3�0a�-���rp��(D�L�!�h��V�� �2Z#��\�w����p�&1�����g�k�0L�tb��s��>y����-���r��)��7<�"���ܣ��l�	�����#�QB�
a�)r��<��$��<�^�1�b"�_�v��:6mI*�I/+�G[ay�E;��Z�A���	�I1�H"����rIQ$qKr�\�C�l!_,!�`!J:J%��u�V�PЊ��R�1�%��$(��nG��	�2M��EO\�a�v;�@�E��쓏���ᤑ>�(L>=9}�y����_�m�>z�_Ul�] :�<�4��/�>�xԬT/�ԂC��r�pR��H��2���9�lW���$���1�u�-Rʌ���Nʇ`Ny���41�O�֗*mݰ4�,���4yFF�[���2��,�)]�r��diI��:�-ߧ���ӽ�s��!;��I���Jc4h=�c|����0������;F���a[<���������y�kσ�b�$�?v"4��B/$�	�������o�.6^.\V�xc�X�� q�`�$��p����ۢ~������J|h
��暖^#%=��J g�N�	"?���w������7\Q����Ld�u�F�-��9�K�� N�'��~:>}������\ϸ����`�_t�X_��z�9�+��Bb;r�di��P|f�vic�.]��V)�6��E,^X:��~�ZE ,%֦A���G[���򳳲����~��,�������"+Z������>_���x5?)�X��Nc�4�:�K�z~g��>��OƧ��}d�+��x׶o������~�E�7� ��� ��>�����(�Y]9]%(GK2���� I��҇,U�W���o������=��`�Ę��\P�г�����#&,��.T@�+��؝�Xۨ#z�q\v��p��^F5OLL޿}x��}�7ݴ��.�F��M��^��c��>N�=]qҊ�xm�r��dV�2m�K�oБwq�H�"��YN����e���6s=��fE��G��B����TVW��j�W~���{��V�qq�ky�����*�>�/����U�<0>u����O���7�e�;�����bK�B�5?|	�'��>A�\nJ���ߵ�/���Z����1 k@-�WO��]o����h���k�oR��׼�����i9�&м�H�~��c�HV\_�ٲ��ıG�X_�C=�c����waZa���{�]��\/������i �W��E웨"=�8̒gql��b̦�e'?&�XY� �$�F�͘�ft�a�}�޶hi�aA�l�K��/g�6+J���7�+�.���dX�ҍ��+V��o4K���/��Gʤ'M��րz� ������i��>_c8����{|�'`�K���X}�
��=���C�������=A1��R������YP����2����?�v�3m���b� ��5`��P^��W��Za���5��2'��_רA���X��������X���k�e���+9��~�<�9T�w�I�Y!p%<7۫mk�@��b@�@l�:ϊ�+Μ)�
Y��d�� H\�X��,�d���b����;��P��ϕ�j3,%���:��n���"#؎ϡ�ٮvg��v��}Čz�����$A��r�����{��W%�da���9?����q����;�w�
�?|p��֮bs=�+{7\����t98���U��;_��}�	hZ�݌)�`����z�׳��<W�)>y�p���e�>EH:&'OK H���q\KhW> ���,.�l�$�Eߓ��'�#��Y���ݖ(ɷ(>@��Y
%T9��D$4���"�5RH�x_4~ܠ,q�L�� T��c��iX/?�+�}?ޱ��܏^�����Ç�@�K.ܹ��u67l�|�o�ƭ?�@��(�$��
1AM�,��UHV*��N8���,�ٴ�D�>���M�oFVrc|��<�\
WN����6T�*:�HY��
+�+u�C�Ijt6Q�`�
������!��휏BwE��\4�}]���agn�F����5��o^w�����g~u���$��w［��QM���o?�[^>�hݑhI��������$H�O��t�5�LT�Y�j�3�g�Ʋ]�܁�@/,V���x�I���D8�4C��>~�G?@�O��nQ�e.+#D�6��9 $1��׺>�\�܁b_7"�[�,3��͞�7T�{t���Ų?z������#8iC3���N޳*Wc���mcs�F���z{6�v3�\��Wi� ���B�Y�*x��S* �E�6�X�S��sj���,�)B'E�"�T@id���A�����B�o3F��	�~H}G
)Nw��^�����w����ci��p/"���v�Q��E��Gd����,��&�̺)[�Q��w�B;@.�۞G���p��g�ueL���{��U������W�ڹ��������S���8�5G
�,x�'	<�L�m @,1~RpP�ߦz�R=�PR��9$�tĎ�D�����f �:׍�{��y�E�EJ���a7CtPOC	�Z�B#	�vWP�@��m��FXm�:>-.��N|<U
���I�v�Q�CSŲxi�,�7y���%. �`�$�g��~�W�ʅg�����N�s��UD5��v��e��B�u�~��x��&�c%O{t�;��K�!F�₇�h/,<7:'��)�s��-�b�� ֖���ѿaZI$E�Ŋd'�-��f�2\$Q�Aι��mX�t�BD,��σ&HjM�&f`�h���*DN
��C�hٌ˹yZ³S�P�m���{Y�,�b��E;DOPEe�N��I�`�G��޺v�0������쵝�b�_��s���C���Ԥ	I]�m�Z/��E��NX������8���y�z��R=%֝�=4Ys-лa-j�,y�ܰ �h�6>�	�j(� ��2����3eH�x���aؚ�g$�(D6-^�U4���rܲh�"�d8l2ta8t؉ _���}���6q�y���!���vװ��*�����1��֠)�u2�I\(Y���Y�)�9��>&e��*�^��M��wX��au�.w���	�TD�r �����ӋHkM]0��%޾�w���(J6�$E!��:Z3q��ʣ/��D�b7��
B�����b�tU��f�nx̥�D��#��w/�k;'~����wm[;r���o�e���s�s�kY�\�7���_�"݄FB!���ȚY���B�b�{	>����k�+[8|Um��X�0�LB]��;��� 'G�����>:�6��C�l^��e����Z(`W�R�D'Q��qe��S�l���8�I�o����CY��#�L�/�o���ɟ.�h���)JI�I�ϟ�u�?��w�$�z���o9|��n���+w�8��n|�o�̓uX�FS�Y,6԰��d�RF&�D����<G�a�E	�ɍ�����]O���Ti�MHԬ�H6��.�j�H��0qcD���]D-Y錕��>����&��������-{7�Զ��x�7J�'&j���p"{`��Q=������>����$?��k�w��n����[����w��_�_{�%��x����b�J�lO:tfW�&� Ȱ���7���Y�f�+1���>P���)�0�
:Nd��
�����A6T>(��F��k��HWh�O�
^�ib`�]#�#���:=�Ȫb"�U�qD�)Q�=-�(�!�����U[Oŉ#��w�<>>u��#��՜v�G~q���;� t|�����&��ǡn;r��n*�2z��kzV�ȭ���/�V�+1��B�*yK뿛�sÕʖ���zv�	tl����>ك�
��Y-�?��}��_�����\�9�$)|�ȳN��v��5O���]���z�U��������    IDAT�⤑n,��'n�:2�/�	+�������;��vp�<P����p�xj�qh8� �1�7-)c%Q1���-E�x���6f�i��w����u1?0E����uo��b�I�Z� �c��O^V�)��.EJ54]!d�?+Nॎ$R�^��KÌ����
Ct#�@PC��c���S���nԀ��&�n>wx��E��~��#>���{z|K������ _w]�6�$d�.�]X#�G.C���tt���8>F�!�(���O�7�����ݴ6R��h2�1��yi�4?|����/�,�T��Z�P<+j��`ua��bqe�$�X��0��z��~�՛��R����9���]d''�O�t��������/�E>�h��q�dj�	�I���nZ<���	I��@�Q�5���2��aE����ܡP����%R%��_���>���d����L�P�ҍ���V[�q�@�u �؟�ŕ%���C���6��#��^�Ԓ݈1�\D�ԣ��������G�&n�>:��U��v���p�<P��!�����YLS�$�r�K?c����fҴ�@1J�$�r7iVc��~�b���(�t"t�(�bʱe3U˓��k���=�+�d�|N��rl�$_��6�՚���V�(��f%9�Rօ%�_z�^�l��o�XIr߲_%�A����g�3O�)k���z���W���xU�_�{����-U�=����5� �^_�ĹY%J8l*Ptd�*���D�DYc������rᔑ
�[�*z(�!a�Bt�!|�|�m��u `<� Q(�<M�;@�GGo�l�� ����L1jSs���4�t�i互����|���e3H0+*s[+f���X\@��\}��q��ARc��_�����3��e��]����E����wrq	x��x�P�樋x��h���RY�%gR���@.���4����C�� �����_	M��-Ӌl�&b�� �t1�<�֍Jx��|�d-m�P��J6Sf�|�-��.���`�<���dE��=�ԕ��3E7�7Ʃ8y��j����Α�/��}�
���;ǼE,��s;%�$ʖ6����$��\�s�I�
��,Ԑ�ug87 ��k!;YҌ�A���<�F������n��t3���f��!�bI����v���)X�fP�s��[�]����Nqq�в�1�Z�
�W��H�1z�D,^=} {�� NY/j�C��M^�ct��1�W>��X|<�d�X�%���U�-*�;��
��8E�|�|C�W��4Q��h3����1J�� >ގ�EZm�51�E�Y�I�Ǳ�մK��m���������i);�͉�4���h���2:*e!�h�"5\��1RZ*����R\�>���s� i჏�M\�}t���[�����D-:Rкs���M0!�YoU�������Q����G�4����1�/le�B�e�Hb�����X94b��J8r��iz����D6�B�l�>>;�P��g�Q���Z.�BH��"�$J��)CYmT���@����b��W����:6q�g8y��]t5[-Th񙫩s[��4����$5XCd�Kȭ0��Ol��g�V[�BNA�{	 u�9F����̧��r�pҚ���x)~S�`Œ�;�B$�s���ag$T���B�j� �Խ��6#�cj�+�3��T�?���q�T����ˀϢ�n�o|V���Q��fk��H0R6��B���%Jј_DTgG�K
��9u(�͵<4 =����WH�պl�$�\�ED��%;�~[K,�sp �����-DY�l�=>%���@�z�}K,���1�lfՊ�\��,���NIb,~���q�H�����&�^�ş}�MG^���{;=��E��7>�!��3#(ԭ�i\f{����T��)�^R�c��[P�<������ۭT�#N�P�AS?�j�α`y6�ŀ��D���a�"	#�T4�(�3���	r��{���sm���5Ց�Y���iT�Q�4�0�쏱�L��>6��=:1{��������]�Wq�i�dq�ʨFbw�0-���,%OK
[M(I��@s`�(&�}����2%q(t�"�6�왢��a'Ķe g�!	5Cfe{;����24�oR�"/'m4�j|O2ef�2<b)\4��cܩDR�5�V֫RU�`=����~���tb��U鎋�+x*�.E5��иg�0���o7V��Igx���$�gmEm3)�� �8���T�<���ֵ����������|��0^�6uM����\]���i�Z��ո�
��jJ�+�
C��'p���;����L>26�g����[��_ݻ��w�����	�Ք=��8���◖�ѿK��p�z����l/�$5|`Z.�9����J�)D���uǌF>�+2��~��{�k�R�G��i�[�.��׬�����1���F]A����j���|6E෍�"�7�W<���	��8��K��I8��N#�/n����g�3��MX��h�S�NE�u�S�j1��GhZi��?S>3�yaV5Z���l�	훹�xC��{h8��Kd�
A+�m�ŋ����j�щ�+�[��?��۶|n��{;}{}�Eמ>/��Ǟ�,�� F�qS[v�w����/��u�P�Bb&�&�⏳
�Q�1�1��)H�i	���%cu�T7��0�Ȍ}����BWcH���3�Fh���7Y��\���z�������-��~������ڪ��+|�((:�����V�c}]a��G�T%;d�#�g�	*3ф�ˮ�����uEIJ��wO���;����C�[jy����/�%	?'[!1'K��e��+�'BSih�n�V��l�V�2��W��͵�>~��Wn_�������8����'�E�O�Wg�MǠ���'s�x�O�9f���@֏V�b�ו��H,[��>Q� �2 �(���]y(�ߣT�P������h��☠�4�k��l�͗-�Q�4�hUZ�u!C|�g�D��NFB|-z�h.�c���R�L#t!�P��g���m�){�����䗶���!�_�؎{���,t]���q��=�A�$���̠\��<R���\o�$'a�FZ[�P���m�m��R�$ś�"
]���r\��X�V�l�'��:svcw��9�/q<+\"��R���'�����+���{
�*!�ӵ���(Z�g��}�^�M)�Ӓ[��^a�UC������>��F�0�0����U��>c����������6*_���������Z=@7�VΊ�@/��N��v�=�w��i.}z�b~|��᧤�Y�O$	�+y{��%�����AZ���/e%Q��������7�k��IZ+@clF�E�u��"JO��pz�(�t!a���(*��s��-ʥ;4��k�}��9
�4@k]����NZ׃y����_{��UB��?���N��XwP��;���g�nX
�Ć�2����1�!"�|_~gI��f�"�%X�B��D��i��vl�@g��}��ss����F��,�V9(4�t�M�j��.#?ЭUk�n8A���H�8GL7~�a�.���N{���!Ǝ�Q����� /
�27��z�d"A%��ZDy�W��������O<66��sF?�2�X
i�����en���ڛ�J�|�y������K�2����Í�$U�a�Aa�N����i-��E>T��O#��9�Z�ck}K�p5ý�$HI��[�j�uE�^65��<��"��%{�x|�4��%R��ؔ�EL�d�NH�a�{���v�p��m,O��Ccb�̢ɶM9Ѐ#�s��BE��k/�0�K\}��8qc/��ӏ�OmU�n���vz�Ɩ���}{�G4�-^�6�jM{�J��A�An�KX�v�`�#���)�����9��X�P�ޥ�a%�<ԣ-WƩ�(q
G#�«�@3@���f�:*5�*���ݢ��)�|�����D��4��	5!��DF@�I��u"�ۉ�����$�c�H���6�t������V��*�c���&���zh�������>�R�x��Pw��a����bRC�-u1\�:�U�O�m䆺E�(�8����V�o�µr�Or�"-^�j�����Z+-�>1UQ�J��rv�k�ʹ�=e䇴��y�2K��� /�f��Y�7���N������B�Q��;F��Gs|�|���6y�d̺c�Nw���5�_����M}Ҋ�������չ���dc}�F���{��8�ht�r�AҊ�劑��j<�8x�"@�j�$�I�)�H�%K�_�R�;���픕�q�R:�b7`/SS@N1�ԙ-��j��Q)����q+�0QJ�)@�O����4�E������]�&z"%�8i�	8W*d��a���I"����k?×.<M|�"���霑�?]�';l�]����^�]?��Z�E
�H
����L���5�*o$�m�\����5�tiDՖP�I�x�j��MBQ��;�hš̕��ؔ�?l0P��J��`W�X8��q��8����xh/6�#�ь�y�br���7g�8훕�8A'�֛p)Z5Ml:�[�����=�Y�i_��8qTz�f{m��s׍��3s���m������[��9|s,B����HK�N=�}�zɪQ�Ғ�dE!d�+�X����;�������]n�t��04�����O�IXb����L]F�e?����(�!.ǿPR�H,e��!F�V%�w|�/�-mAzs�����^�B_mͧ�%g�>޹a@[�����ڶ�����U>�o
�m9A���ڢCaәvY�e��tI�h�aM8�x�T0�+G�HN bU��`}n���K�=Z���	��AϏ�	���T�d���c�l������ul����Ϧ�C6]~�XB*�C�N��]��y��Ws��㔵}h 3M�p������8�s;��+{��E�������6/QJ�ڲ!��4Ѥcnޮt^H��ٕ̍ƒh鸘��O���ZFk/�Ej�Jt�L�u��
��|�">�F��}K!��Q���\��@� r�2�ȬHC*���D��bn�RVc�����q�_Ӈ:0���&o8s��Ớ�o����޾�h[��ڇ_Ľ���o9�4F�腝8�H�7��W K��X�������S�hj���d䕰�S'�2���=��N:e���X
&�43yI:�djǲ��B��e����F�*�� �C&4^�L�$�a���Z}60���_r��;G���_����uC�/Z=�k{��������.Z��G/������v#�+�{��>�X�гe��Xe@�&פ^k�dE�kf���QF��$մ{�>����\����(F���/i�y�\��ܢ{4��BC��^?��^gYe�e�]��P�\�h2�dm�O��3�#�1"��CO���쵫�
��ޗ�ZSs���z	w���	�!����{���ŋ��]u��$�**A�*}#��T�S����Pe\��"�L�XZ|V����5S����T�$�1�����9"��͕�,�5+�bW�� i@�G�BE��l�By/���*�Twv&1�Ϟ���o_�K��'M�ݺv��)������-������i�G	��K�q�[_R�I�d�ܬŝJ2��nK<M��F=�L�)�R��9��y���R�M�>ڵ6D����b�-�Gn1�)^^G1���ސ�pn���[Z܇�>�l���Z����5�u��j�����)Y�/������vM��/��A�c� ^9���m�׏~Z�����-�b�"����������_y�D�G�m2�fhRi��Ġ�d�pF�:����S;D{v��	�<�v�<O�����D�RB[�����3 ��I�����!m���!��i��Fs~QTk��ٙ��h.ɚ��{�WJ��$�O���|1��ZP��|q�Y����Ta0i����p�Eg���Rs=t�����9|ʀ����V,�(~�{/�g_A<�	��1�+$n	���1s�V�.��>�*h���OL��1x�F3�D�>�"S�k��(�Q��;��e#q��a�#,��@�#<_\�k�M��T��~&3��3	�54g���A�=�?Dv����׉�@/���z��Xh�,J�&�>Q�qU�f6�F��J�Y�����>zNڤk���Mݺut��ǘ3��x��}�
]_��K����G0����K���W�0�-�����
6�C}�*��u乙�/��� }QvQ��`]F9��pPЇ`񀀒��iEX84%}�yΣ��f3��p{J(q����C�̦�܄`��ִ�H5d�����WP���7u8-��h��К^��h�hf��-� G�$��Zs��[|��g�#z���<pp궭kW�Gn�m�%�ο��Ɔ�E�W��E���kB�ʕ�ZO�3�G��ʮ�������Qh��ԒuNӈ[2%C�����դ��?ܧ���C�%��Q�5���0,���>��6�������/�fƇL޿55/a���4�m#P1��P(aߌCC��i�.�=� ��S�lJ�BqH��J�bE(5��1�K\������d!d|j�y��h>#���qw�go
t寞�m/D8�A/T�I����\�v�5s��N�@��L�&�w$��3j�@^2@F.2q��/��ŋ��|<��z��伴�ӚɩH�P�a1j]t���G��n�/6dop#����ȩe��`7��w���'Kf��P�>��d���_�-�ZH���Ic�U���J���W?~6޲�"�?~h��UY<�����yO�����|����hs�0{L��19��
�� zr�}ȕK�	ډ$�,rj���tK��� �y�sC��=4�3	��ޞ�JD$��l�^�C���k�Dg�=C�7SsYk!�Y�j�8}<vˊ��v*}}��8&��؎����ٚ�$G$�&�z��4�� ��sl������������n[��9s�]�?��}�9��l��=����-ű#��f�����5M�L��%� �"�3���:�`��Xg��jn���A���Sѕ$�@�1#�v��ڄ
4�#����]��͵��A���b��Q*�y�X��H	��->�p��.
��>ZNֱ�� ��jSJ�z�$�Ճ{�J��ʍYx���/_p޺����GN�ݱv��7W�y[���[�@���y>ր��4���VD	�댏7D����,,p"�4�AZ�!]VI�o��Q���'R�Y�tx�g��2���=b,�SM�0��;�A3�H���e��d_�bY�o�\W||ģ����f
���7f>`��Y.̨.�^O��
��P?{
{���������uU��}�G~n���{}�ȹ�_�����t$$�b�2������K��m��T���:nSgi�&�H\O��RN͊
�+O��4%2�A�]�}@ IL	�cE���8n��%��s>�]\->kl�7D#�M<ʔ](����G���Y��@��s-�����ܴ�A��C�l��	$/>�=[ߏ��t���m�j΁:��[����t�]M�5?|������(F�+��H\�HR�F�(15/VF���J��5i�!��e��LL�bUZ>0� �����-�,T3f�J���KIR+�tƩ����b�jgC�c+�^#��L�'E(3e�����r�B/b�6���$�8�x�h�t�=>6u������8���o���Gp���<����p�=	)��h��1�k
�5�oTs�:͖��pLݙ�&*r87�	�Q�F�ט�25C�q�g6{@,�T��F`'�i� �yF���	=�HOo��)&f�/i��CX٦/4�����C�b�����'�3ߋw��㏏Mݱj�?u���=�{g_��32��9�D�sr���Á�8a��4���Zy�{�h`����7A��+1�(�+Z-��8de���P$Q�)lp��^���t���g����Z���%1��V���F��������z��~P|�)�P/��;)��cw�7:|�C$�� E@����X�ۨ1A��    IDAT�?�}��Ǽ�5E��w��Q�Ƨ�5YJ�t�-���V{fP밺֭3`r��'����0�l�����z���z��̣ٷ�53�eQ���
��Q�1�r�b�������Rd5W���gGHsx�'���i	���غv������z��>o��n�=���������D��Mq3ƅ�0����u��ɨG�9R��2�$'v�Ez�^��MOl����'���������׭?
:rR���x���7K=w&��.S�RN?f4#*8�B�"����������lf�ѫ�5�a���'��p4֡�cwl]�ݺ��ޜ��ʞ�½�xo!�� �!��_1��W���.�I|�X"�M��l�%� ��1�(��S���C�$��A�.ܺ�8��Ӄݤĕϡ̣�I�%��*�M�5a�,�W�h�6] ϭ�("_d�g�i���_�kė��T�Li�H0��2�+�x�1�-�?v����;��ͳ��_�u��}���f��灧5�Ǿs�fq��%e��:� �K�3fz��yչ*���VSB�45#�s��ýb���%$����B�#n[�����!�%��T����g�ϼ�{J}����:ߗZ��&U$)�1�ӉR��2f(kIh�C�:4�%�<RZc��z������p����n���\e^�.|�B��Wc��(-��p�����g]��C���6A*'xp6dBz7�J��Q�Vg�!�d�g�jI�y��j$�䙬�{$J"X���(�fȜK���*Z��I��)�!H��8}�{�$g ���X���b����4=,��#
�R�x����ʏ�fZ��c�n۶f��|C����_���[�.JW��)|}6 ��d^��=Kݔ?�w)��<��ȷ}Ǔi������ؘ�$iZr��#�Z#j�����b�&���	|��$�V�Ǘ�"�sm�Wu��F�|A�9{��2wrzQ��M���L5'��[F��S�=Q:ˉ?z,W��u�i�ᬠ�e�1bի�՜�>�����ܻ}d�n~��{;s��U��x
ߘ	d
_��� �,e��r�J�T��� 7�8E���q
�Z��d�(!�(��K>:Ga��t$�T��|��	�N�9��1=%&P�;P퓬�]#��1�$Opp'JsW�d�B�~
����<i�캗����f�\\�fN	��~���I�B�	�;V��w�oų6�l�/[|ݲ
��if������c`k$� ɔRG&�R������z@2)�2��9< ���$"
���gF3���tA
�&Y�%���a��9Nu�Ke�ų�A4^%y!�AK���NoY��Xd9U"//C�l��]��,ɒ�|%S��w ��ӷ6W-T�|�h�tf���S�T�l�]¡��֣0�����_0���	P̣<�#�V�^'���̢�Ce �V�8r�)ؕ�����\����$�U�W#S;HO8Yz��C\�O��/SV�Tjo�	c�h�`��(����o��M�=o��Μ��� σ�Ǌ,Oē�uŔ#ҳ<�C:���)�$����q��2[�uP���8�\J��q3]<�c7@��/*_�B>0�*��4�����S�$�0}��3���'��$K6���Pr	�ZX
���� ?����-�r5���R��!�Bf̝�2�i��2}��i�����@١�Z#�׌����TRI���J�ТjRO?e�Z��ze��ͬ�U�_�7R��g�S;��p��,ɓ�t�/����XvH~�дZϙd��>g���f�+->^�`2���2IP9+��+C�iخ/C"|j�I�����HL�͛ʁ��3X*��'�-5�|d*c��27U"ې^&�֌�j\Q7�(�7�)X�D�l��?�G�߲s�ȧ;�̀��Α5]o�jh��\ �e��:P5�:.u�j��3=�G�ѥ��GipR+�vMel`fE�cR�a����A�L�1 ����#[�<�㈄!������4��G5݌<`Z����3��s2���ow5b����X3r��I���l�?�f����7gåp����&�Y�V/]��yf���?IT��v���y���3y���e���\9��<O<p��ʨ^s0�t�� ���6���s��j��ތ�s���Ui�&]�K��`��fh	�t.m�+�͢��:�߱�^����׏0�_S���$j�D�����M�k��VL� �<o6!�q4k���-����.�PH����(=1*sUzh�-�c֛FRc�Q�f�p6�X�߫ ������`����߲*�'�۹�.m��of�[��Zrh�Ɲ�%Ç5�eN��6�؛dBM5�%-�Ŋ)�����
d�+�%��˔m��D���5��fX�N_��M\8xv���oK�#p+&uh���R�jVZ�
�=|h���׌>e����f�3s]�����Ȉ��Rms�O�Փ���*���H�2��Jx�<:��X�*�!\��ǰP�]��'���\9����n��t���53�X�}�,�O��(���ȯ$`��*_�q<i��?:>y뎑�������Q���F�_	<3ו�1�V����&�	Y���R���������qI��<8傜�%P1CJ��8Ak�
�}L�3k��Iauw����,.�}FJR'�)����M�t9�\g�<b���vz�g	�YT"!��ue���ܶc5��js}#�Q�-B� z��ށ	<���\۳5�g�!'IY��v`���'x��s:|9�+��n�-�9=4ڰ�-�Б�0�&��ۅ�`�h�i�d0yP�"�N��#�2�\�M	9n_8eD���<�F�Qo�9	��3��m��**Pr���m��r��լ�3�`E�#GXh7�²���ch�YP��*�S��E�*�F�Ɂ�By���qp����#�O���ɢ�!���sJZ$׺�Ҙ,+�U+�E���x��J�8,N�n��EGWE���]dr�7{ ����j޾�W��=2>yێ��ï@m�����Z�w7��\�ç��3!,��`�h3ő�lv��f�1|#*	({a�+u*��l��c9//�8E����e,�w�+���M�"vu�k�"n�B�	�6��2*����@櫨M�ie23VV������C����:�Ǫ̇�7,Mr^�Ö]Mo�`�6��'q9iᵢ&ep���?}���߶��>�;�t_K]�d��'bAx�D��hy��4,��kI�P��FN�4�x�a�4'n��>�'U��̥�^���&7��l�W�H�¤����KB�O/�*��G�%e��&�x�U��ѕc�zB��V����G����<�k����2P�s��Rע�H��'	F��H�>��v�N)I8��j����7n�d��{z=)v���ib��o�3��㚉������yt�Cc({���-7^Hlx����N
��V�{j�la��Dy[T\-҈�e�s���A��43v��G��"���&ȸ��fP���'/CFYO�� �p/
��,�K���˾^��6{��MR�	F?�8���a7Zfc���Swl\�v��o���]�����#�@ߞ��}�u���DN	�h%�/��)�
��3>�����.N4'��Z�.�$�N?;��3��I%))�w�j:��U�ˆH�s����͜ʴ�$�%�9W��㊣�O�k{��	�w��S�)���B��f�k�NF�='�$�_��_%X�XE��Gqն��
�H�?>5u���U4&�O���N��\����s�7YA��0��Q��m�Y�+S���Ŝ=�I���@��c-4G%�`K>��Cȯ��1��X7-����y]�ʕ��	4��S?���?�b%�)����!�BN�z������m8C��˼K9lQϢ������2>Q�;���º�*�>���~o��p��O��y�p��Y\����_r&���v�ѕw��{�|�9쟬��fQsmX��9vC�c(�x���*��/&�x%�[�j��Ko*��8�xo�G&<	ݛ*}
f-D01/.�S�-���V)|=뇤�A�^I"��8��-S����O�M���@����1Cp�(]-�N+֓;2Ά(Tmi0^S�"�ɣ�f�ix�@Y�?pp�έkW�g���n�,�==�{&�p�;�"�%��w~�'H�nx�VvdH�M��9=�v����6�16+� ��"ܡn���h�D?0� �X�e�����w@�U]���U�չխ B$!	0�`26"YHx�a���x<�6�q��	6 � !��Q�PB"�b�s��ʯ^���?�j	{��㿖ׯ�X�T�]}޽瞻�>{�tyF���y�˩F�:D��Nr�f'9S#����,W�����PKr�yȂF��2��]c/WP\��$( 4�k�X�1"2s�v<6�˘X�+�}{kǒ��${f����6kY�W����������$�v4s��q�D��p0�:��ˀ,�d|�x5�8K`��	3� �x�)/b�
.Ei"�R�DR�`l'Ln�&�$�r�:����/�hI��I1�i�T��F�	J@a��0�">���3`���)J����8��H�E�ܳ���
&V��Y�����3j*>wri��6si�*��I(x�]X�2��g"I����]z��ʌ�e�� 
ޤ��?j�Q~M[��Gy*D5�'�)���'�jZS�IG��t�sM"�fn���#��3$�%���r�H�L����#WVӨ<�ϣ 	)݆^�?�c�����>w�N�'�q}G%�-!��Bǉ�ٻ�Ι��k��j[s��[k*>�D��K�!����'~��nzfI��dkެ���X�rV.T@��-+sIGWw���ұ\X��KKW!�ίs3���YA��c�E�$�����Ii�{�!?4jZ�amf��$0�I����x��&@��P��Z繬�OH�A'l![)A7�ZO`�9�y��5�Q����Z�W̬����Wř9ci�-��5��r�f���[���
�")�!���w���4N��s�/�:	�"~�Ԗoa�m��a6�.X��:�{$ʟ�	Wz�B��"�¶��Y-�Zz/�1Dڇ�� p�._�U�^<h�)��K~��b�� �6~�qZ]!��;��t��Y]6|?W����[oYZ*)c�r�Z�6~�n�j��u�̦�x*�iYŎl9;��
Hd���u��f�"u�y�2yi��-�I�b'����Iu�	r�D�{�8��O�5vd)��
"��پ q賯l����#pO�_�Ka�A���އ��<
|��_Q4|�k.l|���ʡ����yz�f�b�F$��@��HdQ7�_���]Ek朻jLپ��z��/��mb��#3|)rU8�$���0g� f���-K��z?�F#{"�h	�?f�閻���hq?i���!89{n��;�r.p��9,9��y�@U��S߽�GV��v{ϲ�V�<4�TC���;��:�U�3﹭��o!&���H��!��?�O�&��R�Q:���`(�xX�iu�<:�/�"�C&�Tb�3�q��Oe�@q;��<����yv�)/��.���=լ^~����%��߀��q%k�� j�$<���YSH9~`{W���
��������V�;��O�~~��Ĥ���*�*��B]3\ΞYr��O�D�E*e� �
���`��>T��E����,�E��W��k�P%�N�H�Y-�5,��� ��?64.��N){���N�d�NN��(��m�5Mώ �CCr�T�Kx�{�������n�Z�������sG��mw=Wfˣ|^��]�?_�Qx��y)������^H\1���e���R� g8�:RLbO�,?]����$�L�� F�������Hw�A4C�� z�a�FI����%QZx�q����^��L��C \���,?'�S[��\�w��R�F��t?��<�_��jKib�WWx�W��v�����G���٫K,�Q�T���7��5��|½���O��b�إ3gm|X20S��%�{hQ��!n�ODX�?$�L*����JKP3���D�,ĉ�	?�{����i����Z��I����8�d�@9���?vB6I�	��hȍ^Cw�<β�K�u/���T�Fm��|�A4TM;L+�������������XU�(�UE�翰?]�{$=!Hf���t��H�&cC ���u7 !7���0T ���\sl�"�1U6�`j4�M�i�0/��@
�
&����R1�}(--A(' �����b14wv�?���菥q��GOt"�r�jA~ L�➁�ϒ��鄡 7J��h��4�t��� I#�v���l^�f��QW��3߿�E���vv.���|���v�����UE�:FQ$���U�����c�gA��f�, )�0�U��4����Gj�d�]�`�8�&��Ȳȿ�@~@��3ǢЯ G�QY^��'���|ι:Ԩ��m����׏�{�E[�� {?8�ma$Ӥ��3/4�Xǵ�&�%�.t��[�ĔJI��,�ȰL�11�,��Дx4��b]�xa����(/��+������;���U��E/lÓ+_����x�F9�](0�5�B�%qYB�ׇ��<t��a�%�[�X<�ϛ��Et�q���2���tz&�>�è��|�8��~n$�M�N�;���M��{��{ch����v�@�x��+QA��!3�S���D��ꚼ�����~�8�H\���0M>����O��cь#>G��ٳ~v����i�c��xv�+ȱ%Tv�*ڃ�x�P�a� ݤ�����{9�8�W��P%bz�h^dIL�/.jn�!
��(j�`�x�d4֔b��1�,̓a���u/�`�M9(�;��J����m�[���f���q�H"��)=:��tD��>�K�?f�={�8�Hi�C5�3�:��Y!�\�ӊ�?�?��Њ��پ���ϓjN�ٜۗ�KR	X�\�K������q=�=Ёq�>� IiV�&�
?SR��	�=!�˯���Z��
a(�/�f�9{t����6d3�Ig4b|c�j�\v*�sY���,�I�3bt^�[��`�e�&�c�G��x��"�����&�&:1�S�h�	�D��ŋ��{ 9$����L�3nCx��Dc)V���p����پ�s��g�=立�9?O�F�}���c���hL�0��8��kECj 9�AnT�⡚���Я�q4P�=�#��t$�!��a:��E� ������W=�;�+/��␂Q����Ӑ��no�4�U5ֆ����+J�����$~��F�ŀ}����N�HG�E$ĭW�O^���s�5H�e^��%M�O�� н9��p3><�L����?����g�W?�_;w����k�ܐ���
e���X�hΈ�qi�A��ߎ�L~;��R��YhX�kqME����x��U�;����'MSQt�9�b��Pٙ����z���@��d�xL8��Dg�&A��x�\�a��4b�q�B�@,�7����(>n����à��V��v����vX��d�H#�x����P����~�^��a&|��v'V�}&�t�:%�^>\�x�,���}Ѭ�ϑj�{f��?���gr-��5�kV���<��#\~�C��o��I��:b5��KhR�T`P+�o	^)�wK�ЙW���fP]-�9h2�C9�J�(j�sq����X1\��I�xZ#�t��uHt�y Cu�>(�4J����������i�~|p��=1l��.l-���G��� �'g2,	�Q��O�#�P��ƫ��`$S��<�{�v�{���<*��gSW5uǶ��.�YQ5���%>r��ge���r/�|�-X�I�(~T_;Hq�roV[�\Ro�V�w��x�����Š�f�(X]$1k&��d^�Dy�_�6���3q��1 ���ܥi1f�.N���+�A��'MQ�mڎ#h�b��}�h�2
dO��P�,E%aI| ��|:��4t)��E�IB�t�,i9�Z���c�DQ%؉(��O?�Gt�    IDAT� j��nlm]2����_N>3���̹sA>�Hiq�so�Յ/��X�5DCov���R�ˁ�`8@B��R�(�e����
�� ���j�i�� :�J��l�zm\2m<
��M�)N���y�5'4U�$	E%!�/Cz0�h^d���o�XO��b�G`�A�,��asS��8�S�۬��;�E�S!_���h;<��jM' �[
'XS	1��W�������o_��`}��[��.}	c)��r�{ZP�D �C�au釈���V���Jl(n���r�zu$\su��m��,��R�0rt�H���btu1�su\s��5����	Tt��B�\V\sL 9+E��M����>�G��}�8�tÔ���[��BmK6Guab���tt�� -�;�
��NY
�z	2�Z�J65�5V<��/~���O�fc[˒ٕ��{�_��S��;�9M����s�ְ֡0�����aL���Iŉ�r��]�������Q��r����'BE|���q|�T�k���t*�j�{�L7ZzW_z!�H�����!����M���T*	�W����ځ�[{�Ic���#�D�R�j~�*x�͵� �)K��bHx�t��`�� Ci��֋a����C|�h4&�
<��> ���e��
���Y2��w�^R �":��6a�җQ`J���i��83܋�X/�f�er�"-+�u`_A9�����*��9B �	CbCu4�z�Y5�I��N�������DYHCCu	Ι0#Ja$|��<�	�'V �yTѐs�$���Mغ��32�i�{G[�5D�!G�BB�F�41�νlJvȎ"������˰tJ��
��̫�����@�I��uj�7��,�U]��a�x
��@��jY�f3�Z�;ƗƣhH�1n���A�Qx��##%�мh
����ǂ%��KS��� � �1~
����FZ6�/�Q?"M��[~Lm&�5^�
��_�7G���y������v�F�ᠹ7��?<���ٛ�(7���5W�&��x�r�7T���t?�p�t/+H%e��"$rj���L�&E����w��H������_v��[8���}y�z��Ek���I��tefU�k��	xYt�h�!!i���pܟ�^_>�RH]@vR�AN�$��Z�p�0»3P3)�0RM\8y<
�2�|*�F��zF�(g�$��m�kWW:��GN`0e#j�غ�#4��T�L�r���rH�"K֒��x��~@�c�Q �����oR�!�+D<T��L[����œ��u4��e��~��i?���!u��ي�V����f�tL�)�2)䲥)�*0m��I�**�t?R�|"�߸��xw��!%k˄��iґ �A�����2�	v:���
��A��T���!�!K"e,����Pk/L=�hFB�v��2m��7WS4g+��(�sI̘���x�B� ̾f��n����ǇLN��#��r`�m�h>6C]���^|?���ںtfU�=�^�7�]p��d��L[��V<�j=%�d��L��qy�#�� ��Ml�Q�Zu��Kj6C�{<O�������בJ%�htm���v*|��=�p��F�"���@!7{�O����{��ЗT1H�O��H�ܣ�L��V�V����(=�\2Z� Cjt��m��6��Nԕh�:�'?�� �b:,5��P�8�� �
�x⻔j�H,/���}�5����;�,͵QO���/lœ��#I+���s�͌ߡj�0��*�V2	�y`$�s����	�6��͈�i�bcUm�w�P?�#hvRr >���($�M�ǫ�.==���6��u!�p0��`*�?��4��hE	h*= i"D�>���S�-�Ũ�qh�P����T?��T|�(͕a��;:��>��>@,M��*tՆ�x����G��S��-�Kg֌�����\#)�K^܆'V�q2�y�=�3��b�@�S��F���u�K�Pa�t�Ɏ���5B�t�2c޲e`DQt+�pO��/��P5����\w#�<t$2*�DR�u���N���HkG�Lһ��K%��cC�����"W6�� �>f&I��k������6�iA:�2������7��v-�QUv���3����]wR��Ʋ����r&bfU�!��CY�Y�B"C @�n���"5=����J[;/'�d2ɿ8�Sx�k,v����SL	$#Q\r�6 �>H�w��#9�03�Zl��~Ժ��Z/g`gҢ�N�^6�@�鄤Cl$����A;��ݜT�ZS&4����Γ@k���	��tl���i����v-�KO�������C+�(���D�rLa>�Y,�ܽ�D��u]p^H����h���s�į�m�Lb�)�qH���ҧ�h��D<ʔjI�7��*��F%j:%R��P�'��OR��N������g�2ԧ�0��F�ݩ"E��ݦ��u���I�>Ē�WBZ*d)w��h���xŋ�W�~�@�����`�~�Gs�X�砖�x6
g�����cW/��Q1��tjJ��;�pn�I�]��6��F� �o,И`s%c%#�T~��4�Y���x<Ν��N2���Q��dS��~`q��i\ɨ� �	�^��!�d*��>=J3�V���a>هB艫���4��f�t��_�*P���O�)��� �p�ڍ[EԡO�Eè����c�2ץ���4�e&Q��#�̓p$���5C���Q���9gO@,҇�`���Q]?�7������Aa~���w�ť�z<�����i�2��-�be��َ�����CQq���}�vs��o�G8�#ǚ�D����S2���+�W�z��7X�=�ë�E��p�OW�O;\ͭ-�Ko]������'�>ˊ����<r�]��)��w�����J�����b�����È%�}�Ty9A�8�zx=�g/Ǝ>��8om|娭�B2a �4�t��H;z��}�fނX7"�}ظq#�:k6��),_�N=�_s!֭{�w�ă}�T���_@�������[nB*����o��o���}۶�@sk&N��@n�ܴ��eMy�@����y~2�5���j�F�X�	�'���H5�r��WkKKǢ���ð�����9�dTS�����d\�
H�&�Hg���1'�T�PԄ���lg������֬aRR�2�3�\�;p >Z���W_}�]w#v�އ��?�gt�h|���xq������_(���1�ՓOB��{�]���U�5�1�v�����w����������)8}T�a��#/7����U�V��ӯǄ���3� bX��5+����W��� �B�b��.l�{���w/��R|����֮�3�?=��O����Ͼma���(*�b
�U\��>Ç�L=Kr���睃�ϙ�m�7���f���c�%�}ƙ�{�9�}��Ť��������͋����k�c�z|��)����(�^^�t4��������K/ƥ�_����!۱�}���z���$)�a�WoBCm-�y�i\u�u8|�0�-^��L��Q��a��u����@,�j�P�I!�sr��;S%%T�L��	�:������v-�u����]�����=\)��̾mQ�X�x*�<>�:��3�>Ьt!��뮺Ey��{������'P6b


�C��{���7�'���Q���ע���D�w��eo}�����|�MX0�)\~ť���EM�������{�{:0�1y�d|�?��s/��\rڎ¾��a���9
�7��ۻ���q�fÛ�F��r�8�d{�T`zJ �AZ	������j��TC����=�N5�%��yЊgr+�f+���̈́�H�0��'����M�p����M\��]`N��#5�[T����KO}�h0�J0�E�j��De%�hm:�ښj�w���dYE-�Z���}H%�P�4��
�����	[�PQQ����G>���q:"ho�nkJ�� �d7��m�ak��x�`zk _� 9�RNr��̖֮E�+�7�[p�o���ϭx��&l\B�k�N;9A�+_�a^Aj@��{�|<@�1�ׂ��|�+��@�t�l$8�v��*(2D��.���"ܪ�E�
�w���&O�����ؖ���d<·h�`L���MAaa>"�8��$<�|H�FgW2
��9��3��������	Ԡ?��O~�:�o�,�g�u�xJ5U*�d�&���t�/�y:6@|0�����X|� 'F2A<��N}4�d"��B����"G��N:�&�T��-���f�1]CV��_K������2�7H��������#�����������M	����4mA�����ԅ'%��2�JF#i��4ɥ�C��)+� ��3�ʆ�N~���o�.ٓ31rM(Dͤ��tF70�'�ʸ�$�(��t<��e���%(��GNA!�f
��툷q1���S!k3A�<Yj���ha�*��/A<Cg3��!\�8����%B����y��r�QS݈|Ұ1�v��� �D�&_2z)d!j�O��Y���kѭ�e�o�p��PB%��lU��(HB��Zw��2L��'X�H�)t?�X�	H�$�� <�X�NB&ȁ�0�fR�$	��=:$_������ 2	�?�N J?'I��3���S> ��Q��I&�}���g�d\v�y4^ȁ��3Ja;2�`!F66"?Ǉ��N�d�!e�P�*!��qU���� 7BNY�m�gT��;|�lނK~p�틋$��|�V�j%��~W@��I4oJ��P���,(�+܅�����<Y�@�,f�L�`ኪä��B�н�B���'��8m�����T$�%i� ^�r4���fRe`�C�Ʀ�(�Dɖ3�%D@�F��kG���=�'�d?s��	"�-�Z~b/�f�&��0j���bj��6�t.�U]>|�U5?�m֒I��մ�|B�&��(�8Xq�y�{���@���a���8ĎC̂_.S�Cq�@�K1y��Nz�0���n���	����C��l�&%���ÌjP�7���׋�^.q�����#���2� ^BFA��PUƞ>������BF�q�7��L.�2����
|C�����3�J�Oh��Ϟ��@��p����?I]�f	}0�VP�9&�pZ�o;�e�Qm���(�w
�2����3��{)�f	�1�:H%8���q�~�4u�z�����*OsӥN"�u��mO�'6Қ'man���G:
Fc��s���Js�+C�`�+���������@�����T�������g�j��5�����G�48M�9$a�����(������NI8���{o��r��uUE��"������)n�I�άf��@T:D�3oY={�q��8m*s�mL�x�`��Q��yzĖ<ȯ��'N�7��M5�D>^߾+���_ ����TC+����{�����3�̞��@���J+��o��u( �́w؃�h���D7d+	6j�UL����J�[��-��\3^�Gs8��p��Q���X&i�U�$!�H��&ġ;�%q\�W��@ ��_�������P%��L���c&NC~a!<4fG�������D�bf�l���H6�<|����/	��f�ZT,���pݎ_����B%�<�e�^�m��q���eF�д�u �]�����L[8}�xL�4	�dc��{���}ba�"�.���`�m����S��������~�m=tX��ш�a��DEPV]W��;yyk^\~���B��l޸	m�\�g��;����h�0݃Q�|��%1��E	�r<�B�W�a:Y������Ɩ��3�?GUs㼅���;�����K��'�L���j �@O
�h��fo �<�k�˖p�]��o�{_�^|�9<��\�~� UلO���(Ws�RQTR�o��8w��H&Sx��G��+��"��RT�Pg�ĂD�� 0U��g��%F�͘�O~�#lٸ���I�8�~��ơ��I0�q'�Az2$i���d�q���)褹��s�̪�{�}s�~��<kΒb	��#O]��&�.Oe���Y
R@�T�lZ�_�Ϝ-:x5*5̸�V�4�$�^�U,�7��J��݄Ly��<C�ct��0B��o�3Μp6ی>���x��o�>���H�)��cu����x�1�(+G,����w����5�����g���#�it��A�џ�D�o�j�Lj���O|�~��-�6�Ψ,��������s�5t�X��6N5�'&sZ(qR)I���P�M���M��Z��'�"����@�[��k���_w-"�v�܎^xA�]:��ayjb��2+�Lh�-�܂q��!��`Ŋxg�.���`dUW\/u�4q�f�j�����7��sgl��Uػw��@�X%]
=y����3� *�m�aD��p�M�L�<�jx�;�3�&d65w,��p�ׇ�N>��G�}Y��Z
ƒ�w�WDhR�H��0펬�H�QE�(uxń�wM�ބ��GJæ�;}q�W��+/g���۷a͚�y���)�p�<97%H���	99A��1c�Hx��9��ˡIkMt�p9�������|yyy�'"X�l�o�F7�h\����q�T�� �(>��B5��4�����A��x�%4�ssKϒ�oo�g�x���S�sǊu�ū�3��Ԉ
M���̴U��N5y���R�3�D�px�z �MJ��_�26���q���!�N��ݻ�v���fɼ�(~�W����<q-I0ԣ������cԨQ����W�a�f�Z�N��;�pW ����lx�/���C����xs��GSk'O+��e�F	�p�D��N`<a2|�[bܓ�zYp�l�O	��WSǓ��斮��-`<�e芝'��?��ʼE������Z��v<�r=�D���N[���ts��آ?��[�b��4@o�G��|E�	=B4���"\q��0�Ha��w�v�KB�%�-�*(,-���@?�<�I��=<��՛o�رc`I
֬{	�w��0ΒL1VFnqR�$���P��2�L��?���b���8����-� 5�P1�k��_6
���;+�قBb�D������Ǿs/��>��Ot.}���ܳ��{\L�3~�3���sV�(���������Ee|��9}�x+�j��٘
�oF�v� �-@2��$\u���/A,m�����ֹKA�� ��J���#�J����AB?�|N�,�Mӧc��q�({~�Kط�����啨��Fdp ��0�;�؍m"�(��ڝ(*�G�/��-~�$�$rN�k,������i�S�qѸ?�i��{�Jl�ib��������-��+��{<���8��gW��Oϟ��]w���W���x�=\E���fdќ�R�Րb�g�T��$R
F��� "�=�y N=gO<[��>ě7����z��_���B�ǻ�:�1�	3�p�e_��Ƒ$��oڌ>:K&����W /��[}]��v�1|�.y1���� ����w`��&8j ��/����zH�"����\��� `��_�bD�?�ԇ'�s�٥>���o��֬�����Q~�Ts��K�������9hPd�����+߄�Tc�؏lk�S&���C��<~�p�	��J�X*��N^3��N�E��:�-G[ڱ����!@�#I^|*y��@~)&$ɝ8!�}L�0EEHdl<r'ڻ!��-��y�H㎘���Q�e�-��ӽ/�6~��z罏�ܗ���ef�1)�S,CsS�]�&=Ĝ`?M>\9W��I�cx�V�ԟ���g��?��{���B��1�\?o�؇g�^V��Q�/q�z�5�=�0\=I�&
�Ɂ'd��ti!iZČw�$��SFz=�OY���$2Z;z��Ð�AL��D����M&���	C�*�� ��^�L�^�  uIDAT>��Ye�oc�;��x2�Pnj��д#���d��M��6Ν|6|d[�q����a*�R�oDc8�HS)�^�t?q�\�p��L�Bbp�~<��P[�G�g�m-=���Ҫ�����ճ�>玅��rV��嫶b��b��?�\6FTI�I��u��G+��[c r��U������,/u�5�t������qÀ�B��`��0�7�`�	>��ilDqq1T�75����Z=�×4jd�Rb�k��&����r��5��q#��.4w� ����cL�ۋ4H�g��	=y�X�K�~͌����iǙue��7�aU��)}2�^����=��_�]՜�ӟ���[f>u^U����p����0�c��\v�&�X��E]*_VË}��$�qѢ�p��A�hif����*T�ֲO���`���	���B&�T���������CM]=�K���Ȍ]�B�=?�7����Ne��-�DG~�p��OG]�(���� �l��(��r�E֫�s�K�5m	>	Q�읱��CV+�m{�{�?��
�?{�6<��~]e�u�]qſUx<�4"�j���kf!��p@� �5����P���v�譔��s �6m���8{�98g�\����8!9���"�1j���ҫ���5�\r	ƌ�Bp�[W���Q,	��٤�����3�$Q���Tח �Ԩ:c����e�Dǆ+�!�_Dӊ �\�-0�$w���6�����7w�}d؁�/����97��|���#u @1Vq'�F�7|W�\��u���(|���ɭ��!��Ǹqg��ɓx��c&�	�P���"�505��,ֺu������.� #G�N�t�/[���O�S	�p�)�V�/���?��5�~%H�α��'���1��q�W4+^!�C������G]�[�����ڿ���|(����?;�_�%��/�{MCI�eye���7�2EQ4K�9Yб%�&�x6�&�7���
rs
���a�	���ۻ�6o���1a�Y8��8�,9ȋ��S��.�5��d&cp���+���'��K.Ec�(�@ze���$IM���H�W�Ds�1��q��ע���TN�8�ٞ�����Gh���(��.;RF�eK�E+Mz�F�2z������ij��|�̏>���3>���~�P@�}~�O$T�qd[-J������d�rlI�=�e�^o�ITN7�.�|f.��e`߮�رu�;�Ǐǹ_,�Ye��a3�B�:�G��!r�q6l؀��f^�W\u%F���(T��C|ށ�h8�r��Lk׮ő#����k�Fe�(�IZ��u����������	(�DB�e[�m�q��X�T��ےi��m*�M�b���jW��������Yvǧ�g�?<���	w~���0�F�?�ߵ�wlg�ʘqc��/^�|\�&JdF
�>���ˤL�������_��e�ې,��
�D�!%]�t��I�����`^v)jG�Q����k�^��7���7�?���Y��o��~X�8n���p��r�����{`��[�v�8��q����m(y�q��Pc[�so���J�(a�ڗq�D4��.8cǎe;R�d�31v#8��i�/M�"�J��G�� <�^z%j+��6��D�<���ol��ށ������I�)�<��w��e?�3P�c�;���6�R,�5q<��w� ,�ՏI����+�u�$��1�7�|���+.Řѣ�LR���8U�<[�@��h<�u�~���~O�~�jT4V�P�����O�Yv����#d����	������2�����ya�>xo�>�ܱ����s�¹��t�J$�&Q)gU����e�A�09�G�����/ĨƑ\��rB��b�8���In��!P$��^y}=�z����W�td%��Ʒu��<�fŽ���&��o}���,�A����م�;�s�7e�dL�:�S�ó��+7H�=��f*8�%$�4֯_�M-�v��RZ�a��������X�� `��߽���(����Z�׏D������u�|�����uW�l��r�/� �㧌���{o�������;�g�N�ȝ:y���ڟ�'2l�Bu:�l��D/��x"�c;t��C�7�4�z�Y��,��q��tlz{������AU���~���h�л����'_y��������?���_��G�
��s�v�ڹ��ϙ8	��Na� e
4�xz��89I�RҀ�믿����u��ѣ�2����)�z��D�<���+/�����TW\}-J�j�tm����#�?�Б���C��M����u���u?���� �n�֭�Q���I�0e�Tq�'�j���� ��.;QHq� ���8~�_I/��"�>v��j�dU9W�=q�_�D���ݝ�C.��
��Z���~���=�����߻b��]��J/�dӑ�m߀w�����O?'��"��k/O��,��e�zަM9Ր���i�0~��npI��!sR;���Y�Q���tu�����MÈ�c�+�㵖����7�?�wQ� �����n�e�Ȑ>-O�v��A���B�yP6�Օ�He�l�N'�f���"�L�%f�����Doo/�����ee\��a�����}��!�U;���ͬ0��c��1oA�z�tN�����>�m��O��5���,���OS���'O���N�A�Ҙ/ͩA��
�S�b�v&�g	���E���2�O���F0�ΐ�r�i�/��B���U�tR�b������Ͼ��}K�_��_3ȟ���f��>c޼�_�Ӊ5UW��z(�J���(Y�v�w�z?QG<�R�G�O���]YÖ,��etH)5��]"쩿�P�վ��N��4��#�۵�Voxs�5����ox��7=�x�	g�:u�iו��Vy-��r��.z�auv�l�!�l�U���h���g>��0*)�D��K�HC+���I�j�͝[7�����ߴ�����߇v�_�I~������^o�#˾"�?�#�!E�Y�H��J�#[��h�#��fڑ,;c*��:��.�V����"����r�$�VlG���H�eiۑ��d�	�J�D���~���ړ�3�V�z��|������������?��C;i�T�    IEND�B`�PK   vb�X��n} � /   images/87fd8349-f00c-446b-9712-cb30a7c611c5.pnglzuP��6�V�(��K��r�)WZ�p?(�-��w
�Z��R
)�����;�_f�L��l���>�$q�����hhhĚ*�hhX+hh�x8�z�gN�UX��:�hhM	ﭰ���=4̽���a�e�5;��hhOO�*����zp�!�ތ�yw�g_\�����0�����(yrZ�O�ͧ�]F��^6|[�D-{����@�RUA@%*ɔ������w���<��kO&�E�U��3o�~�^l��4:��wUp�N�j��Tx��-��)\)�5���Q��V���t�L�=G�霖�lFHU:)�L�ج̐��5	�@�����kV����Dol!����ɰf_��d�Hf��:_m�\�?�3�V�h���n�Ȃ7�{�qZ��$Ŭc�ˏV�S�Q꘵ �&�2"A��Xw@���m� kA��G�eeÑ��vIi�.U��r��",�BGǊr2�~�빕��
�2"���;ˋ��o'EY�I�V���z����h�%ʞ���{".�U��̛� �8s���N�f~�d��Z=7_���K�W讻Rޖ��s��Q%������Y6�����$�]��8��%h$��p#orQ\af ?�M������r<_J���N�����_�����%��j�K�%�'���hF@7^�ğ_����-�jn}��H����)�*�_����h*�|����37������~AwI��"��mծ\O�}�ٛ�j-'�}"�T��nb�2���w�?o�`eϚ
S�9�*c?�2m�P�v���c	��n�3�Yg\��f�\��A�u�\k���Ռ������t�0��_�,�O5iʌ[u�3��?��3��#���Eȝ�A�[�
[Ĕ�K߂<>ͨn--��f�Ep��;:q���ӠD���oe�z����0����H�
��{�6糔m��� �V��81���x�I8��G+%�}�N���Ӝm����������#b�b<cP~��)�����K�x���G 8�%�9Q]�����V��x�E+59�]mj3�ǈ�ޤ)���nN^^��S���뾠����ō��zz�b�m�p�m������:�\u���FD|]�Z������0{
�\A��};�jf�P��s�=?���vQ���3�%��^L͈�+kt}-`���dixv<���6!�x8w�U����Cq}�M��O\��8פ��Im��c\uS%?'4�V��X�z��r�鋺x%-)�ïj���WY�ޭ�Ao�����?����mk���JM�o�f�-��9�z���=[�/� w�+w��g�U:���愜U�T�e���:m����U&�5D{�:l�!�T_S�9� W '�ʳa��>�k�0[`/1���A��VoႱo��]��?��AX>=�f<Y�/<�r��]`�N<|�6o�r������� �|����=|��:Uڸm��[?�sܳ\���v�A�X�!a4v%;%�A`mT|4��="!E��+i'w/�Tޙ�d������Ez��T����X(}�)R�̗�>�0�U ġ�>R5��wXjeqxA~��sU�f#����Ԝ;�QH��a͢���հ��ڬ#�ܓ�\k�5t�lQ���JR��g��ܙ>:I���E�Lx[ז�?���&�[�0�*���ON�W��.j�z����d�rڻ횕�W���j��T���!�j�>���VH�q�;��PeB5�[��)j��4ƕك���}��Mk'Γbm�RV�M*�3 ��Zu�,_�����5�6ǣ&���0�`�5V�/�c�=Y1�jv�E���C�z .+˞�Qr�GE0r8{E�]�%E�h:��xڨ/����s�9�g��N�25����^7JTf�*4�V��?��7=_��0ō�h�O�2����X�����F�I^�q�r�P�PHt�4�i�-�Q�����B���V���b�yyK��@~F�����Tr���=���$����M��ҩ5y���@9=rՙAUN�Ǹ	��@�}����QnP�o?:�p�a#�Q�5>+v2v��p�a�4ݔ&��r�J$�5�,���_�3p}���G�8���F�c��vB�W=~(:݃�5Z9�|IǓ������g��h��:�}ߜ��h�w6] ���K�p�'%ܦ��Ť��M*�̟�Bdg����4A�X#��e�3�, �tQ�:k�ܡ]�|(M����S�"t�} Ks^��=L_���Y����ڥ���H��oN�sQ��mU|C8Ң���a��e�����[?�G��NV����N�u0sU��-,h��S�t���?m�-Cy9�j���W�eH���e��旘��o��{P͹r���g���H�
-�-��L���2s� '����m�����aP57����O>����b�	��[$A�$��|�>cS���d0Z�}�9wf�P�뇎�*2&w���B/��ɯ0��Bq��n+Z��|#�L$��=��d2�ܩ`gY��h�������_>?-����>w.�E�	q�<:��6*C�!�����r<-e���ѫ�E��J�7\���B-���/'i�dn����< Ϳsx��G+�E;�2�j=�����"�[,����2�%#ȃz��*θp|�Vgg�[s�/]��"��AzCL"~v����d�vD�$�Yƽ�C�|�o���r�ki�F�U��o�i$�fo�&��S����sQ+��.��T���1�x�mn&A���n6P�
���,-���{�Ae�]\#'#>-��ul���֊�r?Z��n���tT���K�}:�懷όc�� GӚh��id����� ��6� ¹i�^9=��gb������ҥ�*����{~��"�}��z��td�X@���}
>����a첂�$~*f�
�w�	�JF����߶��R�N�	:X���nݍ\>�~���3���K[u��̔�OJD���:+a|Y�fi��ߵ�yyz�Ԅx��1mi�r���6sW�l܎���k+ �
^|���׌1���ś�8)��P4?��N���CU�ǎ�gi��M�
{.�0Z��>Q��2$������m�ũK���#:���
SS�&��o,K�E^)�	?�u�rE	��H���^���lb*��/�Q��>bg�����^�H6��x�S�J2���?�K��Xȶ9�H�F�˞%:|���z��7���k:�ʉ�%�Ϫ���n�R�I ���Ν����i���&�$w�U���r[�Q�Z|-���t�L�+��c��]7���|���ĲQKխ#�I�k&?j�(�7(K�ء"���ٛ�T�GG��?Aˌx����G!��Mͪ��I8��,Щ�隕H'�85pC�w�淝���@; ���j�ne�n�/Q	���� jv،ϧ'�ڭ5A;6�An��m��Mۥ��hnG���g�/�׭E�D
;с��Ȳ�C#�<�	�T�ai�d�MB	�ґ�Y���2q2�kn*���U`����;d��a�j{�1��37�k��I��(<�\�ʃ$>?�b�ۙR�$vN���ō}��S����$�����O
Չ#�K	��?3�i��퉴|6�Ŀmw[�mʭ�Q�pG{]~]�v4V�н�
�X�O>�,���#�h|㟫��b,������<ݢ�Ռ��M�%��~�KYi��?���e(Џ]Y���*���!L��J~޾� �r�*��7�� �����!$Ʀ��7\��[�E�?\<�@����p�B�dk��D�x!t�'��6�������HګH�a��c�jEJn�)(O�귭��tn�Ŷ<�Ü�4�e�~�1��n���)v������2+��C���}S�O�n��ޞ[�j�a2���,a^g\1J��r��~|�=��]��)�-�C��H�ūmL���mUG������E.�/�E�&��T���"0���0_������� �03Z��DR�G��i�����������'��`@i$>��$'��>�4E�^���xA�Κ�5�#�-G��� �u9mW����c�X������[�:�J�Җb\�Ǆ�>m���GF×���c#[�z�$����@�#0B�a���n�8Ts�p��Я`�.:�nh؜������$���	�Ae�`��=GL"$�� 3��$�aw�;�(�$O�D_]����2�I�ǒg�*�z�a����K��v���k���n�!1#={{e$���hZ�F�I����K���5�T�I��%/VO� FM)#qB`	2��6%���<��gdM�I�'H�ʰW��M��ȿ�`V�h����n~���b��G/m����*܇�<k˚_�0J#_�i׬S��T�ƨ�нO��q��ןZꂓy��=��:~[�h�绱�{�����V�2��d��V���X�Ps�PyCrQ��ji�_+��g+I%���^��+���>]Z��.�`}٦V�OE�c�Q����j����g[N^be09�>�mb�J3�au�vB|�r�Ė�8��oa��X�$-�aX1�A�n��Br���ī��!ʐ�Y��Zq;T��s=h��*���4��<�R��+���m>���V����Y����K���[4s@G Q�|:d^4ST.��`�;�r�U&�Vh:�}�F=]d�so�y�t��ߋ������!�`��s�e�i��^71�w6�w���Ŝ1im�TA�^�_*�'�̱�wH5Z�O!�r���L�i��l��"~��.ϟ��3���]���+I��_�����U�Ru���A��^��x�!?8���������~��j�2��.c?�\��=�I#�-0��T��]��P����v���h�����;�XG9�^xw�圳�����=PL��&�^(�4Ы�«���PMsEi�/\�6�=��P�,[8���aIQs�5����ӖO��`�
;�!
zyOd�G���㪡g_騫*��m�ʧ)N,z��n͡��e�6߹�o Ҫ�g�{�T#QK�,��2ԨR����v#���G�t�Bw&��H�����P��'�%aWz�S��*�hW�=K+��Z(�ř��Z;��ϟV��V*{f-��n���|'��� خ15��K9��_ӌ�'���>%�I���ⳗ��U�?���b>T�p�H!��%� �-���k'j;m�S)БN����=@��nC�w�e�WϧVαP͚v3�����Sc�T]z9E��K�g��&C��`�T;&e�=� "�c�{�nN5L`5����OЬhm��t����#�?�e�fV{'vj��ʌ���(<�;  �Z��(�;��`l�lM��:�|���a7п=�3����g�NL����
/ �:׈�������@�U0*2�|bdx����~0����ek/���j����Q���e���,��L�+�� |x��M��D�bAżO�uN����;3�_G��������v|e�99��q0����U,h�\q�WO����Q.�1Mq앿�`�]�� �`<�K���m��6uNZ�U��bN�U�W�
|�5m�=��R8^��~tHY5Z��.3李��ڽҗIK�O|��e�w)���H���Zq.���(�dN��S(��B�u�P�o�����8��Ѽ��?�X�g�1�t�ֻ������� ����� �ϽT�n�E8�4���8Y�̕��K�Q=�T���anRR
�#Z}�IDt�d�Ig������U�K�JXJBR݃��z���)��s�s�` � Pg�t�;��4="1�����,�x�A�;i̙�"����א�U�f��b��\֮�З�p��I��7{�!���5�Wb
���� ����c �R�=A/����)J�-��F�Y�.�iX��f����xtT��B*�4��`^�R�!)k��ޮ�e*{0A�ʘ�̓����Vy��]�����IIKK6�'<���X�tBBf�{uġQ$~+�
�����(S�7����"��-��Co����7�����E�
q�	��Ms����12QO��N�l�'zo*�|gag���f��V��A�Ƣ���1��*s���Y�K��:-j�"��!yy���6��,$�������O���q�A��G
i�]���A�^����7��w���9�W�?/RǷw�M�yhJ�#2I�鞀RVd'ӄ�u�?��y�RVo��"K��@?ۚ��L�Y���o��F��`rQ�g��;;��1�}�>NBz��nY(%��Ѯ�Q��`fQ�!������u�o�¾�T���7j��Xt��r������ϔz�ѐO���?��噲6g��R�HYvb��2����]����t���E�+����%$���Ͷ�Z8�X��	Gg~D̖�K�S��4fYv7�]�E��NDj����C������׺��+�&p����9�k���~)8���I!�A�g�)�F��S	9�y�L���K
�ȋwP�l�CО�*��,m�cgt�iշ�5��q�&'�<�*��`�B>��<������W���+	���_�{m��Fx�6����UY���z�%�j�ŷ��<\����l~��|�}�]Wu]8B���!�:�p;%����Qw��.�u��^�}�j���m�n`HT%�,���Z|v��p�� XИ����MaD5����mU{\���B��v�z�|~���^��> �r��~o��0��� 7ڰ�W侒�)0	W* �=�P%����U�ߓ�>��;��V9�ĠK�ז��NטVc�8i,�֡��ֻBS��}����j�՝0�.�T�W����»�7ټ��<��3+�M�.@���b�R躟�i������2G/��긋��/����\>��eY�y��Rxs�/W��z�V$�u���mM�1P'��o�f;�$`�H��(SB^��9�V�JjH�5W���d��&L�
�uT���[BEc�(p����x1<d	�/���ץ/��}�0وpz��^b��f	:C�ʳ���nP���f��J�gŗ��D&�|B��Ni�ux>sRIN�"I[]Y�ࢆ)�?wӜ)�����u1
�i�ڪC�P�RxD:�dLY�r�W�Zs�Q��%�r��ZT=__�#ӵRr�����5K9����ݧr��>�\3�N��1�5i�\�>,�����-ylt3��~7�J�����2V� ə�,�=�4Ϩg���c��.��a��%t�L>ju(i�S.��nOʔ5J��MW�ܢ*\���5T�c��+}W����}���(��Zᵼ,�Wo��hֱ0�i���\{�Wxɴ��Ԑ�d��%������I�\'�^���/�Zyu�v5�PXo����k\S��vGk�ak��Ȫ�c�o�O����T�q�b�Cd�����`�����R� 5�[�\Qt^p�<5�e����T�Mf����� �zDb(2���9}{�!}�k�� ��J����N��wb�����ߵ���e���O�>؉���M�p3��8���[��{u�k%9z��mr�����"�KŇ��������gA=�!9�O�ķu�h��>L��h\����[e�o8I�?�	Π_3�m����N�yo�3���㲧o&!��$����$���p������ˀ;�����"�.���)H�j:~^iX�
�tf�c��ey����"����C��Ƕ�Q���{��^�_�]��~^Y<Ï2]�kW��DV1`���-��a���~�]m�������^�8�=\�9�>��"��_wP�����i�3���6�QUh'XaH�+@]�{̲�F�fyݾ���m���jJ3�r�A��]/��o��_�_�7�2�V ��>�L�^g=z�ѭ�o�/�®��+�5N��`��2?��� &wO���Ț��ퟧ;�o�5|G�L0{�r���JMy�*����D��!����{?����8�G�W�R9ԕ�N��0���nK�5������FM��6�,M�m�A�=��:W~��ڹ;>�(?�$,)
�N���1Z��?b�]����n����DHmCn�aaő�����N��9������H�H:��K.�z��O�\~9%f�/�6*��&f
�}ZOGW�d��"k�`W���
E�O��Rz(d
���vIԖ�|O{ި�g� w���7�����-�	E0g	=�1�H������$i����}�����uB�j�Kzux3Iֿ��o�$����瞷�LA9��� �N+�ݓ���8��w�,G���0�1��dá���w�Z;�ݚ�_K/.&�BP�羏��Ֆ5����k�2a����G������&������	��6������0e�.�D�_����;��'p_{:H��w'�*�@U�{�����q�u�? lx`ږ��(=�X����n����xsgܰڸ�m��k�	.)���Wbe�hz�۶�KTE��P����ӌ=ʫ��u��]�Qj�t`�V��/V'�[��f�k7�g�z6�`>Ɯ�K�y���6D�H�] �]%+�+gR��13{֞�t��BC��ɍ��K�5���7݁�ۆ�s��ջ�%�n<�w��ZT�ê�������R���'ؿ���v�T ��8Fg'��f�����Pzݸ�8�}�i�:O��t�S�9%9#M�=I��ۦ��F���*|h9�hy܎W����Έ7�^����oʮt�ԉH�9������h֙xm�Hc��y��.�Sx��Ր�am]��Vδ$��!�O�Dz��:�W�Z[���v�P��:�H�4�*yw�ҠW�;Wc�I�4tn�4�{�.��H"��U>�?�ͫsC?×�ū�ْ$&M������Nѓ�f������%t�Dg҇A�_��o=v���00����<����E��p]mP�eI��əc������G!]�>�?�oa�T����S]�v���E�v� V�j5/������?~�"]"�*g�F�`n��դqn� �K�9'�g�@R��Bg�x"QF[��J��_� �qar�3��5�4���x�sJ������]�	� ?M��:z$����c�dxmq���¼����,���
�(6Ӂ ��%�T�	R�7��j�tӟS|,,O{3}�L�xy#
�ѭ�	,���lr�J��s��$wǎķk7>��wt����n�'���a��*)f6-iC�~�ޞ�]sP� ʁ��E0H1&k�Q�|�#}G��{;��:�;�o%_̉���k6%���.[#��;��;@��Kj1U�5�)b�,���¹��N9L��z'"��Х�S�zl[zR�]�!&����'��N���z��4�� ��R䧷��M���r�C�zq���)7'����6��"�#%*�&�_����Y�NT)�mh����˅7nP���B)��P(�KZ��\���z���/[%��7/,u�2����
B�uY�-�3��1�6�]�;���'�3�R(��p��C��Q�+���U��7���PO:|�l�S�|�"����("�X����-�Ӣ=@pcʈA$���ʤ�R;����4���g�&���&�_��>�(2��4>�He��Xl����uC�zb"��Ƅ��py�D����i�=l�͓��Z2�{$�WP@���"�������0�T֑5O��œ���Nz|�|9�D�;JLM�ܿ�wv̸���y&Ԋ4K�3�F��Q���p���ѽ#qyiZ�	s+��F��-T�_7\�����4���#{IQ�q�&j��8b��0z>���Ba����Ȏyyۦ�Ή�>"������+(#d'?ٶ9B�8|�F�kij���T���/�;�����1!����{�;�~�S�i���b�F��n�_C~���lp��5�Dq�]�[\�7�Q�;�������7o*֊ڳ���8�=]��y-��e�Q���V����d/�en�n�!_H%%d�MkM\�HF8
G�ׯN�����=c$b�#^M����Z<��륄��3�V�Z���1SISo���{%tW��ɶ�zL�W�;�I���꿄�nO18��UL�v���� ]�Ӵ�#6���xXe�~��.h�%�ǯ�V�OB��{ۡC�"��g;t{�2�p#_1�J��W|t!� a,��I��eJ��a�UT�b<���]�o4��**�J��A.��/�z�x����m2�f'�K�JJkZ]u��'K*#��	�L^��;��hۧ��$��J�ʧ� jʬ��ڗ��5���p���}�J2�
���QV��hx���K�7��DW��������奡�a�l,Yڼ�5	�~�(�_��W��)'F02�!l��郞���s��|�3��: Š1�]j���-���N"]Z�X*Qy��N�:����뜖c�/��#�Z�ٷ��R�l�
nx�p��2��g��`zkB����E^|�����G�@)�܏���{L��pjP�.��G���3���AV�=&���������UfD9��j�	���m<f���K�$X�	GQ�}Tf�}�go7ک}(`�{)d�+�D���w?:^�0�#�&A�����o�j�%�S������h�ܠ�1&u呡�z�2���a�{��4#^F���^�Ғ��3.��$�����M��c�#g+s���g\�՘[�b0��r�"�P�fAyh���/X�~L]o&���AMv��-�}��R�]A����\{��7�A�e��IL� ǰ#\}�jH�����g�]�1�k����!��|�j0@���_bZ�0a]���O`�L���B�c??���D4��&��"�Z]&6���o����� /]�{�!�lH��x��3\������bvU��!�������p�vx��ld�Z�o1-US�O_���-"~�ÝF�jL೻�Ј��,���[��"5��U3���)�EI͖�_w�؉S��
ހ�a@.�?��'��� i�C��DD' �r�u[W�=5�Z3���	�_�@��c��Դ��ˢ�B��+N.����oFki���q/]#J�"��~M]B=;�ۼ����R�y[FAA�?�Q=|	/��Ѵ`�E��4��ۮ�'���a���4.f$�	�����!
��&�\!z-0�"�*P�؆f;e%>c��P������U���Y�Q���>6"<�/!�Y߻�E��J��c�NW�����W��j�������'� �e�B�J��bA��3����}��
w�QKv]n�z��Y�vY`�:�=N3lDv-���vj�T2��,�`�������_�F��@�U�����!����#�R�A�&�E�+��R�^(g��}��K-�=<�#8��Nv�2���|��.��8��t�8nqw�ϧ��S���������ثW���6�eҩ��B�Ə$a5��T�OH|I6�ļ�IA�������y˰���:��7�,�ʗ�R��U�}�vMr���'N�'���	��"��L �\���{7Xl���<�:ܦP�3=-�����[�L��	B���U����j��qyE���t�dN)?EZ?6��&���<Sz��0���?ii���ԕ\�l�l���V��>��l5��Ƨ���M���(��Rc��JdG��4|�D�n����@�&��(�;�tAw��2�9y ��=�0囻����`2	��$��x�%��2��x��XU-C̱��̾}"ql)�
A�7��fBз9|�4�1_�j��Í�}tv�!�]*"R}C:*ȶ{������ ��R����6;d`�>Kv=q��jH���O�&�~dvޤ%QP�em��xvQ��s�{ x�C���A5�G���d=Mt�6]����Dl�����dPc�TÒfWH��I[�����}�����	B?����$�m�~�Ca�fЪ����� VH���JՔ<͛��ٟ�z Eq��u���7A�p�|/R�����L�쭱�_��~�T�$�b{ Lv*UYX�u��L��R�� _4���9��Fv����KB���`!1����G[+��~�%?�ȼ��4�b�B��o���*�A���n�<��j'�6Aa�Ea����ˇ}�%9���F8Wb�Dzn@GNu������J��͋$8!U�2�e����YK�,�4�1O�D�u,���&8Mh� ����O������S�o�Ma``��Z�ߍ뗧�-i�O
�ݙZs�����V�}p�H���a���=J�T����HSҰ�Ì�<��?C��O��yZ�!����g�wm�<7��	�!�i�0�
��̥��2m;����9 F����m�ySؓ�fX�L��N���v���c��"�����mUC�jn���L�c�ɰ{ŇT駻�	�y����Iў&tY2�Mh�D|�GMD�8T�ck���)�Hz���w�"5������--o˱�
��Nk����cC'�qMY�7�ހ?�yY3)�W�iH~NG#s����F����|>�9�~,�$�Ђ7�>��f���&i��o,��l��U]��b���[�z����۲d|�&�O��*<�5����N�1�����^�
o�+�����3
��E굻M����D����ff]L�H���_	������G��x�?|��*t]����NG��?����$y+
�+q���s��d�F�r���TP(&�t�d�.��<9A�0I���zNXQMM�;5�dP�r��/5�y��SBR�{�}1_�GDa�f����~QX�����V_5]��v��"��kZ��q%��G�/?,�4���Y������<h��H�F'��� T%sK&�4�xU�v�X�[���$q���O�j>I-�-�@�����q���h0�!y+�8��V��/�Ö�&���ͤ��}�r�	v.�^1�F�U}��{Ѐ	���:O�)���+eZ8��@r 0�P�bc��9v�-�EzDô��,k$�f�r.��1ya$V	��2O9�$G�m»f
տ�t�x���,�`�C�����w%֜i�|n��SB/�Tn�VZ2K6\�Ud
��:ދ��WxS�[��k�zj�-�zj4~<Еt��Zz�g�r\�5�=�Yua�&��i�ix2�@��=i�SK�U	r�)j��i��<�?�>4r}��A���-2�V�tj�{ETB<�6��<���ތ6@.R[�0��	�����������w4���x`�s'��2����Ӎ+o}���[�H�l�:B#N~|�Y���1�E����r���˒�"�#-֏��C&$Z�S��$gr]�.��8&��z(��������Z.��e�"+�K��3�]c��2���*j�P�~3 *k|��r�{tMK�!f/������`��Z�U����Ԕ��XW.Tҩ�äcS�O�#�K�"��UN>
s�\��B_̻���Г�ì�^��ǩͲih�ҥ�o?��w�|�&�P�������Sm
�O�M�
(^�gt:v�|��խl�iq�yП>k�A�Xk��Gn�׉�54�S3u��پ�����N�UC.�g]$�A�2A����٬��u|1�@��p�j�����Q�����G�x����
%E�y��+lx��TE�%b�+����@n��鬻�U޽f�����p�~�.��[��t�5U��t�=�d�����m�1��]o���=�k�U�[��C��lS��j[��e��e:�[D�{Y�>���8E�SDˈ<�/��K��_��vʼ3�5����K���=��4�� ߎ(p�0_֋u�|��<c��Ht$ܺgt��3U4��l	 Eg�(�<�oq��\K܉F粅���'O����p������Y݁-�CR< Ӛ��f�� ��ݪ����̑a�R�8���O[A���f�ք:_�ZeD�n�׎��Q u3�QB�}Y3�'@������C�U�9}o�+�8�=��:����! q�t�k�vD�"�y�RY^��2����R�V�p
9��y�T��q�wu�� #*��sZ���Z���T���H�a��6bn���P�(1�_{����"S�k�̽��$:9��e��`�p5v�k�a���Jao��Z�s����_9���;�5�s٠��f���ཷY� w˺O}��@F%�CkW_������W7�pH�|�:y�\Ϳ�qº<giSE*���=&aR���+�)p0��񑟔n�~�U�G���[�|��-aa&����c�8�럕	`]y��%ƃ����@�{���}lC�S���+d*�'�~�����k�[Պ��R��U:��.���V��@�N|s��kZ0�CN����ϡ}�z@��h)L!�Iٜ��W�g��������f>��L�Io~>�2G��V
���/�/�)�bC�����\ݣ�D�,�]��u�5���g�<R��+	�T��ߥ�sx���V�L�Kkq؉8����R�]t`6�.p�ЧmV��i7K�[�4׏�/���2)�f������x7� x@�C�Ŗ��i0$O������!Klx����?<9�&������"Y�/�/V�.e���7B��:�4-�.��!��e��F@A��K�<�I��߽huh!L�Ч|L��n�%�I.�%Ti��C:3�(���Oen~�%��hU��sZ��0�����E��t=|����HI,X�����+�^�s�jQQ�8쪧.xK��H�:�� =%��юi{! ޢ��J1�S *m�8X�j��b����-�F:m+g�����x�(6�er֚����k9���9g:�t�������������-���Y;:��<G����+i�i�\u�� �t��$�;} �dDΒwg�t��2?hm���M2@ޡJN��pQ��O�$tf���:����t�\�w�5ݩ��@~@�J�4��0�x����l��j�i�9�6��;�NA92�Q� ���g�_Q��Fu��i�^x���:�ʞ��[�[�,[�B(�Ε�#h&�F�/[fս�~-$z\�9�����4�{}���r�D�kL��XN�1�ע�!ɴ���p�/�=&|�{dԅ��r}Ԛ'� ����n���&���o`0-Fۛ�%��S4d�0��q2�S,�	Xx�K}�M�RN�##gۊ
Y�_� "����[���"��$�N6 �V�]���i!�s�YE����f7,���˒��=bhw̎�
=K�	�"�������ˉ����uMp������[�p���~B��>HԸ��[�F� �iWl�IО��ӟ�qP�Qό��Ǫ��1&�v�B�l'"����O첞�u1b΁�[��p1�O�+�Ai|�b��)�I�R[�z�T�v�j���t�,8��J�V����u 'vH����*�H��]�h�X�|�5R�gЕ-�ȃ�� �Y�q+J�L2ݔ��� �C��ص��<���.G���4��q>��6����?��~�2��w$�����K�l
��\hf��I--s���dj	�>׽_���3�\3�0.��7��LPb6P��߆�����V�Ɨ���Zf%W���X��m��G���Z�u� ��׵6f�eF��Y��;VW����w�6�j�.���^�=�G�N�]�����RuqU/w�H�;RL�-δ8~�a����vdI��g;��t�� I@����%���n0��i�z��c���
���rn��6�ʪ)��:T��?�y�E>�����l��:�� �sp�q6� �q�,�ဗj3X�ky���o����4�-EdÂ��C��8�����:�c4*<AzZ�A���a0���f��f���B<�kE�|'4�3�4r27)�9V~�hV��ݫ���`��@��؍2f�M�\6DPE��i��Eή�5��tp��-3+���7�I��6�K�K���k7we���D��n�7���2E�B[��H:���k^��xC��k?;��[�ZU��E<*�T��X��ܪܶ2Θ���|	%�/�^�)�����'��6x��E0����D^�Wo����P�v_�ޏ#�$Z**�!nM��*����n����r^
��[2Ϩ֏1������}͜��^7/�Q&�n/����q�L��U���;�,[�w@����=:�bx� O/6T�򎟿]&˹�ͤ��9P�y,�Y z�����[��$b�yYE�4�����������EV��S!I�l������v8z�\�X,#%[.ɢ�4,D�NK+I5L5�;l�Q��L�h�@��v���S�{5F�zfJa˫ڌM���ϥXho�}G�r%>��Ex���.L���r��M�ZPD����׾-t�s�2K�,7��Ǘ,C�9H)�wvaKY;nN�?�?f�򫎠i���m#���%�;�-8�]6$����;!���7����}��<��Η��k�k����M�Z3MH�(G�6Y��4�l�����2`�%� -7g.k��XTzk��<?���s�)p�Ӂ,��-��)FCP�&�e8r��l'�񬹪(;<'�������3����''�����-�F��X���٤IO�st�FZl���Z]F���w{DG��X��VQ�Ւ���W���BY��zm����=wY��UST��ד�%!LG\ԝ;�\a���cax��dP�@�&gbJ�#BB3�n �>�l��ݩ��������3LfQ�Ġ�ǩ��J��Ls|��v�v#���G��� /ERlsdߘ5�NY�buo�=�f��%�����'F��L8��
�؆���1R#�ިȒ\[� UU��Th�٢a�|��E;ˡt$gtφ�|�	b��k)MZހ�ev��o��4!��g�:��"��<�G�FĆ�0'�El��)�n@I���;4�a8鈉tV�WB�=	'�I��!couE63�������V��JTd�_�H��-s����;�������*Q�)����myl�~�زh��҄8�ĜA����E�hf�%�3jT����9V�g�=e��Iw�Ik1-�܉�?EX�Y-0/ ��L�G� �-J:�3�>zu�����v0�`]��
_�ZW3���3Xq��"ۑ��Di���iL��o|���M���a�S�དྷ�he�č(����.B̫n�W���ܒ��7��eYaã����nA����3<�ݷ_=��24	D%���	t֕�s`�6H�D=�!u���� �����Uq�@2�`�'�	̠�9a>�'��&�RQ���d�1Eݾ���&Ö1���"Z��Q�d�@QL���%�o�������B0pTdYU]�݌ȅ�C��󫜪�"}�4�3�}z�s[��d���8T�|��z��"�%��J�FF3uT	Hݻ���mkW!q.$��"~����0qᢡ�ّ�R%OPD[�.)�/t\�����֡ǐXuj��>@+ϔPX���7����A��+QG��$W�=�.�����AuO-��D��%)La��=2vW)� �̖J-߆{���JTg	��k\��s�c�5/�("�N��d�/Z�݊�g���$v��W�A�Z�hS�?Ɲ����O�
x3���D�`�7&/9[���?$��w�������NMG&��ׇ�x;����:��Hp>q+�m�M����i���I2�3��j�&d��M�Y���|tI�u�1z�P�/`��~rK\*YG7A�C4�`���f�)��:yB��K�I���֥i��0�E))�R7��/����:�U�&�x���K3�Ȅ99d����H�<����Я�W����ڦ?r��v�.⚒J�/�IL��U�j��W}'A�1(����$.A��dty6�
O�'���#T�8cؗ��}����q�G��������'E��Q:�Uz�8��h�*�[��尔�,�(���}mO���w��J#"��ky�|�G;����lpq��*�U��|]p���{���l�n�&�D��~Q��3D���<{>��S�5�P����8Ƥ�&#9��HF��9G�Xe�%?>@V{e rnY������MeU���1�ϏS���E�Q`�� �� 4,�.%�=�N��;��M���=�wU/BLk�s��(�� '��b�,�5��K�����C��3�1�`��1ޤ��N�Ӽ쁣���YjP�pNr/�8��S� �n����i�9�.?�9�_/�:]:F�jhsR�'���:KF��zjitU����@a�̹�C4�n��ulې%Pz��T��Z� P�6\%ԤO�T5�&��{>�`�O��cª�hu���u��"�DX'?ڻ�H��o񎖽!�ܡBg����C
ol3Ƭ*��PX��?A$�o-�m��#�D���n<o9�`�-H��:|A�?`1J���N�c��,���:����*�%�Gc7��t{�C����k)��n�������f#P�A���Y@��<��_��!ũ��d����OfH7�$~WBi���Y�+'I��V���{�xH��v�P��nڱ:2�� yV.���T:�_'ߊ �b�c��ֱ�w���j�Һ���gt���M�~�~��KCa��%��&�X�27�1���~g�ƪ_5��[�)���]x���$g3i��}9�[��&#�����G����o\W[d0��i�J?R_RJ �/[-��H�SK�O�M���8��$�?G�K�i�4� V�Kg�[����E���
�N�PS�9Æϰaɒ{[	���=~�wF.���#��8#�:#=	��H-��.w�gn�=ee��n;�<f�$���������9JW�D�v@�h�O�E�߿�vY��{�cTd�{cϼ��<�R�*/���wG7����yz%��T�%��u�T���3�&=���Ӝr-�"7Z���X{;$>����Z''��1h��.�˶^U��f��s�4;7�)��Ծ������Y}Jz4t�}�)�"�Fr��g�-j�%#��+N���c9�-�d�>l�"�~t��XD����t�7V�)����f�E�UO,g=�<:r�K(�� �O�a!�6~���w���gS�i�.e��v����:�N�&����Yk�"����6P�]��1b����Xr����iw����:ʵ�X��=�l�XR�������bK���*H��KG:�(�qT\���h`=1�;я����z{�@��h�;r��bH��.ed�8
UpXA$ d��:*{�7�.�M��^2Bu���˃��?�:��/^'?'�P'�is6nݨ�pg�{�*�o�a��Qe�.F�����u�?�!�&�d�����o8~}�T�A�}�{��.�9��e�K?Y�����BJ�g::d.�ޙ�~9yxW��?�̔�G��Ie����VU�#���.q�]�;BDQ;ac�/8�P�|?��� �vOO�ɹ���,�J�Xow
v��)$�����~�/�}"��h_T�"m� �����'RȄ��'�����H .�������zP��j��Q-�
��ٱ��*�>^)? �m�8b���;����G�U?�	�x�4۟d��J�)���ɲ������S�\�,�㼕P�����"�Xr���0"�6jN�y�K'O<�@!Џ����H�c�䱎��o��M��-�;E-�1����s[ˢΓ��f�a�Ρ�u�h��4dX�ѿ��ŬE�I2A�Iǹ�~G�k��z���̿��yt7Ԩ�q�=�(�o�3���0m�-�G��,~RF�8�VoӜ�	ZJ��I��JOA��:LG~�T�j��θ��"��qI�QI�0�O1hOmOC�*���)|���%� 4��P4�3Z x`�{�ss$���r&>0P�(�8
�ŕwQ7F�C��?�y�
�/��Z�"�Z6}>��wv�u���l�Y�e<���Y��ɲ6�H��9����2D�|���C��G���J�h8T�|�K�i�M4�n�ʀ$�Sh�G���l8.���\b���e�O�@���+��67߂b�m��Y�y��H�4'��)"n��wV�4
���� l,R�N�>�k�
RbE� ]��@��R��}�e|c�hզ	)�<%�������%`�}vw�P~��g|�?�*;3�Z0B�E�7���S?��a#�?<�F��yQ�� 淎����q�l D�g�fi�J�ƃ-#�K�����@p�ҡ]��՘w�H�΅P����/���� �
`�������<Gڰ��~�X	��ؑE_Q\I�B�(�F�����>O낲ժ�<�
�o�?b�"��C�-p���R�d?.���$rc��V'�d�|xVR���ȉ��̂/����ָ�Cb���gCPQԓ�نQ��۸�����a�?t�F�3�7b����Kp���v)1�J�T���O܈JE�P/�t/��7�cf���1�|����t�15�;���҈e�9>�e���������g\�u*��A�l�Gu�C9^:6g���/4)�g��ܕ��0����c��B�y�v�v����.�3-����+]q����[@�~��4S۬@�k[g���2n.�k���/��8jE:507 �.{�K����X��&K�E?�����y_�L��PTo��MAʫS?�����C:T���'xIc㜇^�9��dVb�3��� �n�>ɭ��R��`�O"r}_//�
������@/bź�����g���E�Wq˞�LT�2U���iT��G�>�9P<'�Ҍ�Dǆ�ģ��u4���l��E9��A5�f�9X=.�������M�~��L!qc3��=���l���XI�B
�8qZ��߽B���b�l��)`,�5;���2�_���EGt�v%p�U��:Z�T*��>��o����_0Pg$������e�}�`��AW���Uԗ#�WX�J�ye��g�*!��猱�\��Z�f�ϻ�"�a��!G�ɤ��l���aK?�S`�	O�&#a�ѕ�?p�{���̓&,��ک��n�?n�1�� ���;��ՓvMb�w!�ô?�`̏�[V���r���*����1\֟z�a ��Oa �v�ҍʜZg�u��֤Ц3Vi�#�?Ze-()��Bb�f�1{}��G�Sf��k�gZ�L?�]����j��?��I>@�<�I��U�2�.�݌�-�t����C�R�6�0N��㚂��`��f������f�\���\�gH���; ;6�,ճ�7�Lk�+\�y	��a�M�X�`��S��4�{�~�di|�Nb鞿�UX��1����E�����l�D���F[- ���0�+�|!
�bt��Sxپ�"�F����k��Q��c=&�#P���B��g�5?��2� ��e�^��4$���8x��#��K{���
Hx�u��c�u��3�m�#�����m
*w*���b"�l�#)��g]�Q��-?[��OtW���iX��aS�]�'���J���z��.��, ��zָ��Yؔ�2ʔ4�-���% �`xC�J���a\fn�ws0���L�5	?�����n��Z Y��A���������8_���9p� -	s�޴uQH�*�ոCn���aDy"�̄Ȏ�Phj���\L�]�7���t���"�yWQB����-�y╫,|�`}��Jx���rd�tC�%���"ZYݴ�������s�6v��91i�yN*�u�zw=���U�hQ��C��b��[�k7�����y�AI�~��aߨE�F�8� m��v�?�	!g�c辴T������
��#+���e� ¤'Z���Fq� �E��h����'��A�V������xn���D���L�e�j�2�D��S.fk@!�W�KA��GՖ-�}Hxs�� +�ڳ
�-������~8�_����*0L�[py0��A\+.���͏�c`6����h�T�����.�{i+���G�O�|J9����|������]�ui�c�Y'ih.�`!�MD>� ��Q7�V�ooHI}�t+�*��7���1�\�q_a<�:��\5�Hp��v̽h��>�6G��y�Y�J>���m��Ƙg]����$�/�D�*
\�7�����.�;ŌqGC�i ��v</��ɱk�w"m�n���w�k�!�G��)��?	l�[���	Zr.H��ɚ���P��_8��L��|s`��-��摾j��}�N]p�5�tMGKe;�E<�A�q%)
���6���|��Ye]tk��)w���=�ai��Ӝ�'��)~�γ�« ���{�����"�!ɠ�������g��Ւ����{�䝡�=��E,*:���!82/�V����-`tW%�͍7�N��7]祑W��~��'D~6!k��x��*s�=�����[@x��M`
�݆o�v*�ëk�c�}ss�  O�Y��I����d����$�(��p��շJ�����N���5g���]���X6�We�n��gTU�:K�[������
�K��:�ɼ�/-qd�y��1��B)^�����V�5%��OJ�ci�'��A��
`�;CVR�C�ց�4�����4���<7���&�s#8a{����5F�c��90��>�-�p�|*�
��hG��B=�W�l���o�+݊��`h&��W�U�|'&�<5�pw���?���T�N��@�?�ZDF�'/%2T%?}���c��ƌ��3�*��]��˕�S�����iz:��a�8��R�V�Zej�F�� :�K�C�u��)��Q����(��x_e���&h���R�K��bI���|�2�@���}�-5KO���c*�e9Ek|wQp���ci�����_���%gw2F�ê�w؏(��0��]���b_W�����Ql�/ru��7�r��I���O!k�6!���&+��z-��/$��ϝ����m�����J��������}��\@�ބ����ҙW�l�QW����؈m|���K�`��WXbk�+���=��x���w��M,=Ԝ�N�����ϫ�I��ze6>4�m	����zd���S������/�LiwZZTP�2�K�$A�OmQ��4����3�8��A��}�(ʚJ��@4�|&� ^���2�{�9�����,iE�4S�
��>�C�����4됍��>\��N�ǀ�%�*����,R��E}DIL#��=��J�x��c����L~�d�G�
Yݟ&�M)��~�N��)�X\<Z�4wc�M�����b�)�u�tX����X���wˊ׋бBQm�|��tV�%��5��2��ܰʗ�aۿgdY��:�'�X��-��\�DCg��<�l�DI��j�E�4����I��Z����,�v>�ߴ/\zD�&"Pޟ�TTS8/�\�8�����+���)����n9�.��>oM�$d��v�^h����S�U,J���XɉoЦ�n��E���e�/k����7'"+�f���f�dkU���XKi��L�qt�[����v�Jp�k�J]�=݈�tPv����Jx^a@�.`�E�|�e��Cv��Jtb6D���c�BY6^�0�E5��f]�Øy�v݁�V]�2�%��M�sd샘�
=�ý�\wk�+�����8�ʐ������zU��Ȱ�`Dm��i�Mf�qL�4�ˮj�����)���\��QX�o(W���_�O&���|�Zb l_�z�>-���6�츛XH��"Wn�����=��Ѽ�
���hͩ�0��8Z�?�$Is����WjA�u.��}\;�6�Tx�����F/�$F�������U��ٶ��~8h}�j�Z�H�ˌ��e8��6-� �L^ry7�Gᯭ��YL�	!<m�m�*3��1�ַ�G/D]���u⒲��������0`(�ë��W�+H�1��g����+��w��(.4����2ݸ��<�7Ԁ�]���E�^GE6�<[l'���R��-ը �"d��X�q�ޟ]��֙{4�V4봚e]>��7/(��<�w�_}�?�N�Zp���¥!�+z�x��H�R�궠�^ͺ���Z�y� �P��g��10_�=w_��NO�V�,�?�4f�X��`5������#h��V�ߦ�B>�{�v�|X��Z^�/��z�~������	�ׄ�~�����
���0us/I��|fQ�q�k�fQ��cikE/4-S��ߒS;�B������%�&�q�;�4��+�y���{��S8�꣮漓��?�s�uB��	!#޿��6Ԅ��G��:]�&wX�j����v�n�-�������p��8�Z9D���_��"�����.�ss�m4~G+T�~��� ��j�VE~b�ۼ�3�u3Q}�-4`��oӶ���>4�F�bb�����Ǽ�z��}���j-|�箂����B��[�{ڠ�]y�z������������&k\���cf+6�_o�(�����4�H�A��	��T��a%;ls�'W���R��d�M�t���Ы�`�1�`�@���=:�.�|�1��H�%�X�,r�)Փ/�y̦0+�'��0s�~~,�qN'� w���9c�����]���[?�U�8�4�Ǔ�rK�9��X��e?�eӺb�F6O��/0�!�t�ͱ��s��x���R�5���������%��(����.@�v�r��W���=\����3���N"@����ӕ/�qϓe+Dx\V!���_w
�6*��ч��O4V���_#Wj�։Fc~���1h9K�]~j�����[�s���-�,ş�.q���S��^y�G�a�3/K	Fk����z1LIBI�c	��|�H��56h�]�`��P*�{é�<����Ԫpo	_9yϵI�xըz`�\%D��:oř��J� �2��/�%���'�q`R�|XO�i<��J�H�w���-���պ�d��]{[n�m�K/��;��fw�.�g��Ƅɤ��5�4���Z����$�˪a4 ���@��X�u�U���ƨ�۪�2���7���un��pp8��-<��$h}���0���O�GeϮ+�P�,������QF�Y�8Fݪ|&q���3
>{�_jMJ��$��ߺt���Ez��]B��:�[�K7�QTÍ� )&��=�̩P�mJ'����ͦK��ؑ8G=o���#���q+3�?�5H�z��є*�F?�G�{��y��y����V��K;H�.�zDE(�6��H�� ��mk�(��y����:}��u���3a�"����[剞��VY��}"�������;+F�\�-n�����d�>� �(!�7y$�d}�@�pqD�1E���x���vy����b������� U��>��5=����!�{]�y���f/��T���߰���@�����w������9�'T5���J<�f�]���������uk*��\�Jx|7�q��[)'��iV	�~Oy�F�b�)I4��Du5��Y;���i�S�e�X(�q�"�("T�&�X�
r�
��{>P��^��l�4
�8��)��p�3"p��`�X3����A���/NŮ�3v�X��Z�I�b*�؀�.*�(��LY"]�+<`��V�{��@�ą�8��a����i�����������7k� �Fbp=/����x�cK Z�B�Pk�s�E�m�.����G���SA�՗!���n���KC��(YÉ+�6��m������bxF�&�q�lפ)t�"5�$	��{vF)�ߗe_�Z&�4�ts���� j��{�@�C*y�^xb�T
M���__��h�w<��c�E�m�4��5ȇ�Ծ� ���<_4xڲ��Y�4ᏫM#*;
��okJ�;��=�]a� ���+�"���Nv$��OU #}�
�bu�7LnH_#f7*CH�ݚ��:���a�+���1/�If-�P���Pb�v+;U�z�՞Nf��.��cӻ�ʊ�=X?�d�µ���	@,Es�?���F�[%����+ ���ץ^����wd�5@�������`�--�0DY�s��uړ=��Dyid��m=��\G0?ݵ&Б����x@�Sh���U�?l���Q��Yc	9/�Z�BG�zhND��>����~����=S���&��ܬ6$��n!�&M�N_��T�NKq����ŭu-�a��m��hs< ��I�W
�kI�Q�&L�p\~�O=s ƞ�I� �?ޮ�E��%κ�-���Qņ����OL$|�D{bW�ȹy�"ƿᓙOjԼ���+qm�P��0��Vn\���x���|��O���^�-S�����Bf�X+�rV���$}�˰6�8~��nX�C��(��Us
�n�}�f��Ey�<����:�5���D�8�GJ�u�`q$/ƭ�(x�tn@�?)�24$^�o���>gxU��%_&.+�󬿳�T�EEӪ(M��L
�^Mu�
����ے�!te=S�z�&t=��f���mL�u�%�ͤ1#�!/ҵ��1����o�ڵ�w��Y^�b/�Mg�_U_�^`�*����<���I�)�,wd���Ѹ	�h��4hTb��>f+�����PO���ͤzcZ�zX�~�[��j|ߎ���!a����R%Z=��^��$!��PM�ZL�����A�G��W�t��w.���m���H�P�:�Ɍ�Z�+<�%���vG8,��H�/�#!Ԑ�)����6>�֫��FqqS	��J����s/#~h!M�x�\C������:��t�k�˸ʢ����{�ڥJș�9*�k�w��c���j���iI�H��B뫀�J�Lhkɨ����������j=�G���ӧºB�}b�2����DG�Kc���^�1��b�Fb+%eOk�yh��`�Ϊx�7�C�8��:��C�cu}���I���Y�^w,5͒��	�� �Ks�����on�At��;�FO�W�/��XC0�fR�"K����:3U�x���T���Y�]{�_!�=f��Z��n���1�٘EyMh�Y�g��8�a�|��q�-�t�5#$�/W��=��	�����`�0��]���)�[�����AoL���׽<�D� "��6ƺw	D�N�,kd�f�@LǶ���+�m��Ț.�����t[�rC���}��m����Z��#��MR��7S1f�ҸԺh$��K��lh(�x�^i:%ƺV��83s�Gr�^)[F)�8���Y�]�<M'��-�`:Sa�}���5���=+i�Yux�θn��K�v.jJ���Y��uK��&�Q���~��>�5�|���&(O�C��c���Ƞ���򯥤����d��'��0��1���ym�iT���7�K<� E;(>�s8�n��H\A�҉��@2���+�^I�������d�M����4�]U6���Ng�{����qh=�y�q~k;�ڕ�v2HlhN2H�Q��D�V��D���m	O��J%�$>�e:��+�L�:�Wgd,�R Y�?L�k`쩋��sw/�"ո�M:ԕ~-R8Y�t�}��������Q� ƿ�d���V��;���܂������n΀�N�b]^V�x$9�Ff�Kܚ����^���09���Ǜ��ZI=�dkJ��(ވ��N_��b��?%D�@���({lO�7���V7�~$f؀_�a<=��yF�g��Ϳ"��8��t���?�m%�\����U�m��_kפ�Ǘ�ǴNغ>?��L�(�0kW�%eV�qb�ɿDEw9��E��^W��k��a��L���pk?�]}<X|F��85଺Q�=�`�(�`ı���RX�i�m�p���o(P�f�n�H�|i^$����c�?ϲ�����1i�k]�������*��������_i�l��&�/�|����/A�?_:5���u�݁���P�� ��B~m��#�Q�|��yȟ�5
���@�g�����de>�"_w43�~�0?�E�Ld�S�q����|�Z�����l��`����ow:a*��Ы���eI��u�ɕ�=�=4v�}�b"�ݰ��DG�z{�M8&��A	6�g�� �Lmϊ���5��������2$Ȏ0�������\���إ��L�J���(��oյo�M�l�*QF0��]zߤ�I(�[�����WX�ȓ��wLl3���(��7%8�� U��h��旼�8�y�N�vLq����
����%.���H�G�vieAh=����_���\�������h>�"��X�A{ dy�&��Q�"��Zm�n�� ��2��I�%d�V�]`S���J9�1UZ������;.>��R��C�	{���4�X�0~���]W�{��E�-`�.ɚ�l���";`��÷�L{*�U������lJBn1Z��_�uJ���j34�Z���_�0���d1Ǆ�����B��I[�Ս�a�Z ��� �?�~H��Ƨ�K},�>���L��;��l6�=�З&���Am���d��s�8ĩU��sP!wG`a׈WϞ0PqCV��u؍� �����%�{[��/"B����BDg��Ii������>��{����zc5 ���/�;4F�a(���?X���y ��_c{(�l�^'�^aw�M:����ʋ"�~f���j}zn�L��i��Hg��Μ�\�&�BA/�*�5[��M�w-��v�G�#mX�.Bw��Z)RJD�]�[;?�[8ަ����ɶi>����w���ݤ0t�{s��T���+z��C�O�Y��
��P�|ۤ퓸���ǫ�3�h�n/s��m���Y��ح���N�iw��u�,�q���/����	6RP���ڴ���w{�����Y&���N%}%�AIߴ](N\�9M+���K�/UE�vR������D�)��Δ�%������U�Q�lvinXׇ�g�[6Rx%�&T[��'�l���j1K?��--1? �|0M�W{���ؽ�F�����n�q�x��礈A9���gESv,C"a0˅J�y�bn�TQ<��*�x3OKw�,��]j���v��hw89j�K�=�g�C��z��ǉ��2�+a�d3d��~��_7^7�Ex��; �5�T>��YU]�!G��WU�;�Z��� ��Z�·|��H�q,N\�2���� �AO�O�O��6��~Vݔ5�?����,�J���xjes�Dp��K��Q�N�����ق�v�>"��]^=�dGm��X201D�����e�۔:(�A�!+��+���wD�`xy��P�WRV�S���:��^!�\�+�~,%m)|�?��Pk�av�:�9󻿡q�#H�����ѡp�^�M��Y�AX�����>t�>��ޕ��	��mO{�$=���4����s�.���~�}�W��Хms?r�Du>ِ�%a�aR�EUu����&���I���-~�o��$
y�!�Ƌ8Ȕ�-����ʜۧ�+6�ɨԫ�]@�.i݅C�:�3W��ʈr="�FP���X�,�>� ��৘���J���f�W��;���*�t~nUs�F�O�YK�Kő�� �7�*��sҐ��h�B�}�
TLӈ1�Z��&��q��3,���h�?�u�Վf^hQ��E�
��y�v��U(���>�A~����e@r+���6G,,��AXQ� ���ɷp+6��+��4h�]�bW�iH��fXk�-�b�#hQ���B��k��q�T�*�?��,j^�,~������wGE�Y�}Ĩz����(�V��_�-�?O�q#V�zޱ��|}+�~��X��u�u�9�,Z |m��v�B('�Y��nو(Bg43
�[�R8��pUьJ�i������k�˓�x}/ķi�������l�>�L���p���q��H����������w�ݙʯw0o��*.�Ƌ#�E�YzښN7O�6U)��7ހ��N��{-?�u���.����$[E���̊:��qN.P'�s8%��N7k�<��Wu �I��	��|���K��[�{!�J����C+�kڀ{�踼���kF���F���o[B5/����`����U=�=�S���H�XQE�5�>��<�&yQp+���I���֯rj�'�|WxN�I2��p��+R_߁�Ɯ��]J*w��Vp��'�?:�FH�q�
��T���bxw<�=�-T�b85��ߙ.�Q[�Mz�r�$mћ'=�*�BB&����%���:�D>�ZO�σ-�*1�y�<��q�X{�a�Y]��ܛw�qJ�iP�j�Q,dۘXy�*	v��8Q�^��:�mYmM8�X������X�Ƀ>*����z�-�Ϝ�t�:���@T,�"<z���29���#Jf��ӿxk�g"z�ڃ,�Q��~t�|o��:����-�'��ő#6C�5��2(�e#��(�����5փΘ�+a��G�=7��A�K�ͭ �7�A_�|�t���xs!��AXC�$,��t�|���kJ �D�i�5Gc��մRz�Ϳ�������H{Y�]|��Nso0���������|ᵊ�6)�8��Y���^'3� 	��"m�ح���k�+"4?��"��X��f*g>_�%�P
T*���WZqV/޼���!��̠����/�W�$�.�R�������u�b�M�����}H/҂|��W)N�R̅�2���a�?�d�i���5+�ޝ=�8��w�"��N�E� �(\B���h��'G�Y�^���G�wӆԈ����;��R_\�Z�:���������y�<�AF̝�cA􏝆v�a��ip�f��#��{��\�f8��OPW�G2K��A�=&KI�|/���R��%�pY�F��'�R>s��%��Y/:���ϡ�9;*�m-}D�O���TVf���U8.��R�~��-�j�B�.�.]�=������*�q�*�ԡ'��(mD�_[ǃ�s���c�m�e�.R��s�<�����B���P�����F��I�<�O&~��_f(��g�2�)c�@�GS�Mp�[h�x���DB�{��͕��z����/_�:IX�<;�$�[��e��p�8[�Ul�"湗}:-�7�v�*�+j�'�#g^CV�o흏jU��,�n�?�7�^�k ͙�Kv�SOčS�H�j^��E�;��U%n�A�E��Uk��z�%^i���k� /�s�ټ�[I�@�8�6-�^I���A���Әչ��)5{)�xq�e�,���5���3�Bq�6	�[��S�m9ϐɤM\v�f�g9X��ti��Q�A����ʠ�zԗ�:�3d�.Ś.��XI�8�v@U�ހ��b(��+�oL��V\��!�M�����M�m	o�dh�1�A�*3���/|#O����ײ�&"�Q��`�D�o���K�]��6��z������Ց��@~��Z�>�����er���	��'��6�d���V����K<|���	��_ط���S��9d��RL�ZfU76WMΨ��lb'<n9��<h����.i �M&KP`m{Y���M<�,������rib�m��&�b���U�j�|�"64�� ,��o��$��k�������
�[>[�.C����ďp�<&�r&!ήk��5%��T��!sK��U;����iToF�r�T�W-�0�����7��������+���=��;�������2�A���B���J��1V�KX��D)�B� ��Mת�HR�K��I�t}���V��@"��(��T7�)63ا�)��2 ��y�<.@�:��t���k��P�Z���s�u�k��I~�dɉ6���M'��rZ�Jl�FB��$Xw�e�!wR�(:�=Ո�t�}�;a<4$~�\
gR���<��[���58j�C��d��j�x�(M�J6V+��P"q����u��K@����b߸E
dH2��!��˸;6���i+`���Am��_VFO(>���F�]�9�)G
�l͝�B�0�C�F�A�6�v`P���6=k��z��m-?\ղu3���yyd��-��Zx��͓əO XQ�L^P�~������]���i��y� Z����W*.`g4�R�y�x�%�_$X�f͊�1-u��@���(ߛ2�R��|Kq����������fn��aw�9��6K����=�Y����Ʉ�l�暋� v����x U��B�D�@u�|$j��L|����8�=�H��[G��z��l}c��,ԯy�{D`7%ֶ=��d��XHwn�b��^��� �@E��h���WC�o�ʊ�4���+��Zrc����ˉ�{���h,�.�<zr���^�R�y���<{��%�ш������6
��Z=����6�c����:�_ߙp["rC�?�]K������3�"#��SHc�$p�cL��-����#���`B.��i9�>��{���j}�~�I������b/�}�ڵcZ��iR�'q֙j����|�]�uL�H��o�.��2��<��r�A�S�� �@s���I�r�Z������6[����w���`��2q7���	J'0ӝ"�`z�!����A�]�]$%����Ҥ�_��(�`��Ad����!t��hD7l�*s՜J.��k�{s��u#`"ījĮ"#߷�"�J��%��Ƚ�F���p��� ��}�Ӓ���4ŔA�U���������n1׻�0dǄ�ǵH6����Z9N����#�FP���l8�Q/l"����J�:�V�b$���5]~��k��_�^��iu�vy����ϫf��p&�Y�7�k-L�2D,��Kp����辪��;m��E1 Mm	dW ���6�D�Q�gE� �u����ב�I��	#�5�[
}�Y��~��G�7���=oo�ƍ�ƶ�ƶ�4v��mۍ6�m��m��>������^��9�gp��9�&�Sǹ��z�q��v�Í��폙���	GǖΉ	��r\�U��N���%D����u�%]6���L�������I��b�&��9���|;ܿM�ܾ���$�M�7�f���F$����M)3T�=kn�(�D$����#�ݺ��Mbح��H
�r�+�q��4���U��w��q5����֛�&��,���G�GI��"G����o�U2��;~�l��:l-���>S)���g��k��͍J՝�Yx-5o6<'��ko�p�GE�I�M�n{Fm6�}";
+U4%'0݅���mZ��'Y�̅�����.��n{x*��MxB�t~�V_��a$Ig9A������0��oW�o)�U��S~舠g�'�eW3kX#)~<o���O���٨�0Vt웩ƻs^P��B@�S����Ӂ����XP��8�uE��¥jIkQ������{I��JxR�q6��D��Y#�~�kj�Fh��Rsb;O\M�˟G��u��<-"�_H�6��&;��� JL�qc�
�Lⵖ��Ex�:�w,�3�N4#]-�ex%���ا�J��@c%Yy<�VUN�q�<�N~�렿�Nq����i�'~���� ��/�n���:U/p�띫�\[[��X�����D�\����I�4��o�����xzgɧh�&o������z3������3��k��e�|H[�zH+G=�q[si�wv~��10YE�b��-�!����������`�#��V|T[�<���R��m4�A=�Q������d]��/��0��g��Sj���^��T���7�`7R�^�&y�c�Q�6��ܾO��tֆ�!J�J�$LuqS�J2DMX�G��H�@jA$	��d�^2�iV�n[���V�|�I�h�i���ݗ��軄*�Ϙ@��DE���9^�b�ƩOɞ|%U�W�Q�����[�93�(p�^#��&�].:%Qѵ<X�o_�����a;IB7���
Gn�y�~��aŖ}�ٕ�f'�=6Fe�q��u�KR�޴;���j�l�9u@�[��з��N�:�8�[P�U.�e-�C05�Z4�X ݉W��ЇW�����61O��aS�a���QE{�iň�r��]����\�����,�My���8��ݧ}+Z�I�ӆ;؍Z]�6o�^ߛ�Rd�CYlb%dƵG�Z��fd�	q4:�79%|}� @��RϖٜG7]��QM��t	3@A��O�3��"�Ί�⎡B�:�A���ٮ+��M�����C���.���7޲Q<�=��E�a���*C�1:mu%3�s�ei#���o�rv�ϑئ�nyh���)hJ
�h��/�*⼝o{����,I�l��Uh0#'qx�ֱ�(ґ~�l�z�����,�Ԉ�3�?��*�^?�V�m崛�բ(�h:��Y���bK��4�ҩX@*�m�Nr跈1_S!|��A�(�D�������Yרi�O�_��V�J|��*$��շOG1�
n���Hɴm*;��`����^E���p�>���
��]���[sY�I�H�e�~b�
|s~�)���[�z�|��s�[k'B˳h��d~vr;�����ں.��D���-·r�%���a�iz,6�~Ts*f��Й �N7]�7D��A�
j�3U젅�}��gT�w�_7���6���!K3[��<47����w/�*�
[Ex���槝��ʮx���A�D�G�:�^c�kqj�����
�r�[E�����)�����N�����C�)��P�������THޙ^��(�]SM��o�`�ױ�~��s觕*�d_P�*⊨Rm���J�:�i8^6�	�*��M��t��V��""^JE_Иq�A��C~�Qv\1+��^0���3��E��u&|�Q�r��8�Gk���"�v��l�<�w�G�y#�Ő8�H�/#��x���Vd<�Qz��6y�2��,y�Ȓ�Ik�s�t�M��u��4��x'@'F����{���/]�l����^PlR\��P����-�wu���\�e������mRA�c"7�{����E_f���]�*���=7�/�%�@�[���AWXI�!���ǼA9 !���,Q���Vw(��c���?���r�>��m���pk�bF���D�-����&uh�d6��#���[�)h��~͍����ῇ�]�-҂�Dڪ�&R�|�%][`�.?����q�G��e�y�n��FEt=a�q�Ƀ�;)e �#����`3�QgK��f�ۖB ��K�3� �?7$�t;L[����[��n��&�&lf>H]c
�=��OMwMm�TC��=�-[➖�~�P8�����%�h�7k�>B�i��]_e�� :"Zn�a���$/�'z�V��%<\���h��-��~xE��(5�,5�f���x��ZQ���n(�~�H�5]�]���c��P��u�DTlRcμ�G�M\c�&r�,�'��]�pD���t>���/���U�0�lf���E�.7yy�_��Z�7�y.y��\�6Kx���*՟_���FaDv����P�[H}�~د�W/��v�i�s�>W{���l$:�8~�XK/���˫t�`��z���m��<ۦ�?z(���濛MI�]M�����)�z�iX��*�r�i�`����!Jt����dA���&ҤA�I��h�fcTPV�5M�Μ�QhIM�}��;ӌ�BѿB�;�>�6��h����jԻvKk�1�xJ�j�G������+=�+��͢V�Ʊ�EQm0D�յxNJ���`[rhp�^��I��D�⸒��ı:�k"Hݯ�t�����g�Pr����2�x��168�Ir*Sy)���T�/��6`z�*QX*<Z��Z4�C6��f�n�nl6_e��(��)8"â�����L�U�n-�?��n�A] 	tA��V�U%։ۯ�T9ؔ���
�Dy�sm�5��V�/vi�䁊�C���	���c5u#�������AQ膷c��4RaNqQK[��V��Ǿ������א@����3���<��w�`��+L!|�f�=U�"��\�������[M����)�e���wp;��45��
�|�ĩ����p��XX�� ����'����1�c2�9�Np�;
��
A/C�M�!�r=����ü����߆bmU�^x[�T4�cƺ�>A9�K���Gi����e�,���UP����@����LX���(��ԡs�׸y���̜�����K��Ѥ�*�������5.����L������nA�/���(�}��aoDN����g^��0�<���?�=tja�:e�+����8���8�ӡ	�Ot����6��W	O=wO'+�׮�����d����{���'�F���B�/�� 1�G�I�7u3lƙA}����A��ë��/hp
��{l�i�]������ �CE��\]��F�}�Q�y����g?%)��֐�.Q��P�
u�Qk'�*~Q\`���<3�7Ȃb9�J�K�e@(RV͖�8J��V�炇e-���C[���P0G�ϓ�}��G��>�q��4\sQ�d�H�n#�;���gl����-/�������(9�ɽ1| �I_�糲-d�j�D8���(�Iӭ�'�������ߑh�����= %an%p�6X�L	O�z�p��������T��7��)�0��nG6X�"W��o�e1Y��u��&C��/F�Z��ż<�+�MRl<�4�����:|������S,���?6�=��wȞn�����`�ԈF��b�2�m���5K'�{����{v-�?�"��E��Diq��C�3��������G�.�9sF���7[���2�K�m'p��iA&	�A�݅u3/���ԭ��Oh���ZdFQڗ�g;�1�t΀9�T���<�X�j��/ᖽd�K+k��֔xB	��}L��[6��
��#�`�J�rvj����}�����lg�+5��)��h	g��� �p�iS�H���#�F�u�_ ��[�)q1A=Hzv���[�L�K��*����a�Y�+9*T�,p�0�	�����d<�����`��/��AT���`^��K��/u�#tݾw%3K�a>[)��/�������Buc?�5:��$zH�HU����]��S��9Y�Y���5ʮ�9@�ZU�\��q�[�|�hG�bGA|"���Ȇ��m�|tcz�Z��Z1�yb0Q����-W��,�[�^�ܛ}���?�C�,��:��*Dn,:��N��﫟ZD�b0�֖;�_-��D�4�e&|��8�����Qb0yZ�,��Uzt�F
y���Q���Ϭ��eʱ(�X�.�?M��U���|��s����PΌ�,��&m�p;W���;��L�$����#�rvG�Ö{��F�#\�ؿC]���"J*�ۭl�����^��[-Yt���2��%"H�iW*���	m'�S���3��c���`~z�h
�z"i�wq3΄�e���t�A^�fȯ�x�8x�@��(�)G�{l�#BVy{a��Ļ���d�#�]��}��e+��A��6]�{�������<���@@���k�DB��[��㱢����D�2��,�G#��u]%��5}B��ۋ}X�as�r�A�OD�	��aK�-�b���U<4�4���ȷ;��b��c�y�+�����p;�ت[.<H��~tʓZ�xn�`	8�<{}u�}^W�	�9*�e]���[H
���,�t�#k�N6�*��8���!R�
�(�vb��ti��?��9��q_���f9]��8���n!��l-�k0���Qoj�6�&d�DTȧ`��;��Mh�.Ct-|C++'K�Ÿ�[G����>�ؠ���އ��[r6j���z�֛�N?u��oCf�yė�,ē;�G�qI#bX*�1,H�.V�*���f���pb��F���Hn�d�W9dr�;*����\�ia����t��@�V	w�h	"�| m�y]L<���<	E\Ğ�ܐ�zC	#G����U�YlI�u�I�`bOPM�ə$G0_�+jё�g!̓�5éނIO�@����Q��:��Pq�!�a(��pI�O���|�t��JI�g�I�,k�(�[vK��� ���:���l��~�����v����͍u5���^���g��M�ܪ3>�q�t�^C5�<C�|.o�ͽ�N�쬈?��{�d}j����q�r�Ic@F�~���ݷ`�o�-QsŜ3j�X�{��;��Ol���|��t|��A���"�oT�`w�s�ɺ��P9ñH��|2����P>�d]�ٚc�ۻp���������7.wi�#&̖�wT?�5�}Wݢcׂ� ��"�������`Q`�).�R��kޗ�ˬ+�����W�aǼ(�{C�0[�B��7��?�'ա���� Տk���ބQ#��^�>��+���q�?���qB�s���{b��L�C�m�I���&���]�&��"Y��{1����ϧ�J)r� �RJK �QVe��N��+TV��V���1%�T�����ҊXB�|����?���ѽR����>}s���1�5ٌ����9���U�PH�t-r^dp�?��h��T�6�2�i-�$�D8RC^ޑ�|�C�E1Q��D���!@(�2��/d(����#L5%J�#�1�u�4���TZ�F
��MD?[jI�o-�5r*Y�\uu�
���sli/��cy�q�!O��.��$ ���ˮ���D`�wm�Fm�Sm�)C��ƶ"N�w��%C�C�NN�ٓ��`����ovc�����̸|�t?>{!�L{~h�����@"��Jh?��Du>>����΅�^���e:R��5G�`Ͽ�D%��H���8�޴��~��5�����
�BO�Q��e`��*�����AD�=8�!�I��5�3�$�Bc�,1:Bn��}_7���EC,G�\��wj��lP���h�~��i+uf\�L��>��A23�F��i%�Ǔ�Dr���X�V,Pg���$�ե�s���H�����L��d���^�����壵��L�nyY���QS�3.9��?l��I���k0���?��}o���Y�(���>X�w�A�����I�EHB�0�l�Xl�2�H�����x��mU)o��
��U^��*�j?���y�HO�M�s���j"�Ε��2a���Wp��yPUw}x,7�x\ϰd��)�ٝ��sG�/ͬѢ���T��[�z�7���	bw��{��4��#�_0]�Z��LW����,�̈"�݆R<��'ȟ�=���5�w�c���܄c���R?��`����ɹ���Y��*���J����7���aJb��@M�@��O�_�2�(*ʫ�!�����CCuM�����!6�����h��ҞK��#����������.m܏�Tp��jw��iJ��GF9��O��H\>�$ ��g]C.Vw���(0�0�:�����p�/|��O�:fX��)���r�m���P'��I�M�/��E@���y�`ţ���d�Ҭ��Y^L�s�¥[����¬Gժh���^HR�V�^-K�c�&&�OpT��2��AvƠ��,����������t,���s���F%;拙��7|GDP�_E>�*�D�΅S��v �>'y�|�ki�X��v/|SO<[E��m���p(S����=}��1έד���"����h���#���$ՇO�����(�rL���ȕ{/XyQ���b@[�팹j�#{�\�lP�i��2^��U�W����x	�Ĝ���6����)�M:�-�I�����3�&��0\��c�0�m���'N��lΈ�ճ�y�,<����ȹ�0�M7x��8" �z�����0�F�.�a���^|��c�o��c��3
��`��)���e�������7���6Uzʟ��mH�0����Ny���XD�*a�� �YJ83ͅ1ٍ�ʐ��(��
<&I��Ҡ3pӿ��`U_�%p7~.�������# �#KwlX��9w�R�F�$e���gǸMۨr�Y)��A�a�ں y|MpJZ��_���]���nF�
���jt�_��w�L7����`"����J��e�䈻!��ʡE�#:	�TU
u��yX�� �ŀ���vD�r_�\F�Ǫ�Q�J؎E
<��K�%�C��j(y��M3NХk�r�8_�M���T^�,a�/�5Y�!�w�͸_���%�(���*E�r��o~��m7	�g�iH\s#�U�nQ�Z?EA���f
��`Q#SqkcKfk`|/�%������?N	ӊ��u�3:ɛӥA91g#:���Q�'	�ܭ���
 �'��G�C��-��(��Ԃh���t��݋��=����������8���L��ߊrI:�c4�o�'km�.�M˘����ܽ����a-��5Q��cz���k�GN�	��O"���U���������n�L��?9̅�YzdM�Q�����p}|R�z���
&`�Ƭ�y;���E
��I��%�=0��n��[]� ���=���MP�Ñ $a�	�����ܕ4��u8���ϑ�{+� �+vUg���-�-i�+�p�Ϋps��9�ͱ�2P�$�Ʀ���ܪdQ��O��*�9����"�OM��qb<��³H�0,`Cj��ۄ�z��e6�.L�ѼԻ}�<y�6���+��nl쨬���$�:���������5�NhF
�B�V;$�7]�a5��\���[��&)��K��e���֯�iy���"�j��nc�Mfd�MC����d����f2�����H!�	BF#�s��ϩG����W�ʤ��[������C����t���WU�������)�S\́����%Y �Q�����@ȕˆƲ�U���R)ۢz����Wț痟d�7M�B����q�s‮*�mI@�%턋x8�'��TQǓ���P���p���OT�U���'��pZ!0|P*��p^ݱ'���'.��X��3��Sd!z�u�h����p]�M���@�rGe��Z�����ij(�0
I�1F�@��E4�"F��6�}
�Ά�c�9+;Ƶg7j��$��b�[.�*H���A���zh4�-,6��Y���u;,vs������\Mw΁!�������>���A�!�7��M�͒��`�S�m��[�Q�����P����;�V�A�?�.b�#���z\c�!���eW�A�R��F�RP%e3ѕW��d/�zz��ڌ[��5��.+�5��g2(\V�ۧUcPs�ňTZ�K�ۘh&ϭ	_Q��{^$&�(��"�?��/fWc?2E\ړ.�1?ǅ�r\΋w���r��j~�M}�}�!H�AΟ��/FW���ᵗ�k�yn�=���݇Е/ϱ�
@_<��ܭ)�5��!�IK�[���|�!z��&��g2�D^>YcP�ZN`-���.�q~�D�#`ћ��h��B!j;M&�G)WI�S�u��?�
�QզhM��4~wE3��yN�Oru%[@��;���@�G��jii��0���n�v��J�Y>�QF���;�h}.�Ö7D��[�q�0��%񜸓���§�ѝe��V��(�wC{�A]D��DW��ũg��
m^����~���Է48�Y�Mj�e˴a��fI���j��sS1q��/�������~��h-:�D��c���;��d�.��_rD#	��
ߗ|m�Y����.56ǘߙq�n��	{� F�qi�d5�81ߤt���<���W_[�7@���=�)���_���L�f�	���
��w��s�r����u�����X~���r�����_Э������+��@���ϙ��>#7q�"�-�Z��v��<~�D�>/v��)<~;"�dC$�j�d��`������ً�Ȁ�GL��ߞ��w�6!&��힝��V�Ǎ/ͫ��lC��w��8F%��{'{ō���lRM�=~cW��Ҙa�\6\ȓ��?�^�ƕj˜̡ }�>'�o����$҉m�����9ؑ�W�����*0:��=�F��� d[�2ԩ�t�16���;� ��Ң&�F��7g�3�&A�!�7b���m&5J�	��;QϮ+�L�:�q4��/�x9�~�Cc[o���7R:��O]ϸx>oY�	�LCcc�{0�i�ka�(�����n����Fz�8ƽ< �^G�X�œ�j��V���V��)��V=6G���_�H��K�����0�X�N*��5�����;~�2���Iv[
���Z
$�d(v�h;��&�)��]��	� E	����S�&7OIUκ�y&�� u]1�c� �!>Ή�旲���Ņ��&�k�I[e-L@�W��Jq��u�W���y�`����� {�c��vv�\�z��z��(�;68<8F�xh��t��Ƨv��C5�C(7V�3�Cx	h��V�u!6�������L����gj�vM��W�͔ڂ`��֔�)9����͝:����Cs�Wl�~��#��s����8�V[��5�C�fvSQ.4�~^m��	t�����(����<
�a�4 ng|�/�Η���[d���Q����i!br������X1�ڥ�?�bnV4����]ш�4���	�[q�F���u�w�y��K�J��U�JL�<U��1#'�V��8�/B��9�< ~�H������!���g�p�g��x���~���g�*5�,� �F�>���g�TF���/=�D�{��:���q%C��0i�Rr����<iV�?b/qww�pea�n�]��u�=W�]�eӆm�<��HU^�8��
��N��"I��J�ʣRA�5ڭm��!gl�N���#��W�V�QW���<o�$�&��3j���,�m;�=diH�	�4=t�|�����MQ�)�����E(���m�C�~M��:a%]*��X�G�g����gG"��3=�D =�F����:xj^E�]�#�6��{���c��d2_؎��r����5���fO����&ǉ3Wu�C@\��@��G��L��Q;���)��։�� \�pYj��=\�j-� ����t(u��@���\���@_�����71e��l��S)��(_�]FE��~�gj���F�W���t~��Fd�wO�L���M+�*	����z��T�RR")���G����T��3>�	�o!�Y

y�l˂A��}��E�j�_����6��{���/����De�S��E�o���Z*x����0���u��,Q��;��}
2=���ńt�(�5�2p�Y�$)~�hy߄��@"X���mO�����Y��/P�N0`�x�U�����WFހ	G�o$��pRҾ��'f���j������c���7*Ԩ�m���C2o�?�>O�%���d��T�ʒ4�U'�������[ɀ0���9�a����K5����U(BZS��`l[ٲ�n1���8>���??th�z3�B"�����;̢ӗ#�2�{��>�ЯE�/��Q�u#�{��C{/oc�9�&���+n��MT�ٗ���5a�U�H��#�������J�5����o�݉��W,�1�rqa��{�/�z,vj�r�[��#Eۄl�W�f�����D�P͂j��Re��1������+hh"�j^�ҽ�v�����Ãs�;�_���T5��@I{fpp v"�b~J�h�T9|8aR���/ST�c���� ʦ�h���p��;��3O�qM��ew
��`~h����{��)0.��ũRW��7���U�~M[U�CmT!�>������Y��	�!�R�ب�v��65h���5j��\���ʣ��A������t%�ޥ������������w���2�q��?����(�L�?G҅����M�O�'�F�6�%xS�׮1����r'u�H�� ���vZe`5� �B�(�B�bRԉ|�߹�fg��o�9ͅB3/�?j���������]�9��|I[��c�`�	�5k�;�����I�0�9�@��0���c�W��d|�f����P���Q"���Z���1� h>��"�7U����l���4��o��OG��hyPI�C����ۘ|�ވ������p�2�$卍Nq6�G8ŘY)t���~���%��B�}�oA��_=��c�_m����/Խ�{��O�[��Ic.Y�)���}
*6b��p>H����3���M?�����b��*��b-x�S��4��e�Jɔ�+K�BC�M����#Ui+�Gߋ��G��!��=y�g�"2�"����ҳ������C�u�FPA;˩���LV��~_<I1Q���TG�ƻ��T{�N�t�[�ro�`��0�DU��C��@���(���(�⛩-D��e	5M!_��D��-I.��Yn�<�5����s�-+A\�,,�:��&;O5�O/�=l!��[Xni!N���KAڄ�׬)�تv�֔.&WSo�yS~�J�GHho���/࣭%;�X�>�׻S���I�c3����im����lB&�*��p�/g�|��Zk@o>������8n�W�L������3X��#�1P�r���c�N¦[�u�W�W!�O���d��w�q}��y��/��/��u�zT�����_=���=Y"�5���5��xǸXo3�
]O�G��#��[�q������'Wt �����x�Mt���>,���>G��

�-9x��jr|��?@��5�<�*�r�c+K��f�!��Ҫ�iז
�g���jr��}��a��l��h@�t�i>�s��*�6Ϡ�$��dqʃH��U��a)w�@ci�>^]��A�\�kû�o>������7�[�.�8-�aH^�����[��,է��0��Y��o�jeEYq��eC&�m�b�}IP,ZOj�K����Ǭ��}w�B ��z;�*ϔ���.�%��̄U�&�M��*4�o(�vS�lzèv`�w��fX�^Y�6�Q�f�)�3T:T�لA��W�d�^keI鯛f<�����w��?��
�3��c~��M�u�:�����v/mF��)q1$�Da��4+:�q�x��䳵n��W��Ӟ=��E��?ݱ��1�@"�P��v�p��l/Mn!�z3=k����Uh�9�J��UI����jG�Gן�6��&�d��\��C�.���|QPq-t` k�G[��d� ��"���#�dM�K�M��j{Iʊd
���Ǹ>��!��v�d���81�@�ۙ�iZ�|�W>eK��sn���e�5��(�g �,�������\E� ��Y;���-u��ŀ1{φإŪ��5>�+��R�I9��R���2p<�V`6E��E"nx l:��kᄷ��Ae��� ZW�����~��8��L�?6Gk�X� ��ù�1/����)��>wb��t�8Y�N#�2֟hNx@ �]ķ�u�D�k^���A27��bռ�y�s�^����?����;�u%Ȫ����m�����M���Y��� �.J�'4X�cb�� �c��9�m ������k4#;E@?Iy�g�.��
�ڔjce�:��{p��̱�����#}q�NN>��N4�]t����"�Y��g�ٕ֓����Q4���3����6F�i�a��@���ru>\G,��.I�,}�F/��'Z��c;�c��E�g���1v�g�:;=Cg��:�שZL���uU�/C�������(������J��)L8�D^ܱ�0% �B~sZ��}1�a1Z�/ w(�5�S���W_�}r2Ė�=���.
�<�����X��2�*�$�uL!�%��d�Y�f����;y��mqQ�����W�Ԓ�9w�F��vsٺk�j	�ѩ���15�H#��������� ��L߂���9��~���P��|��Rcl� *?��$,w��|���w�Ɖ�l���]6��$���S%5al�=�޳S����`1�V����
}�Fԓu���î���x�S�-�z���29��O��'�l�&iK��@����Q���gb�X*�b��&k��[4L�'s�&�Φ��jS:Qr&�A�(A}y��֝�I����������գ��LS]������٘Y�&vm�����Յl���`4ǔs�[yu\�}�J�����J£��'o��4�o�q������P2tlF���@���L�Y�#�u��	`��Vwqz,��{�����j�f�P1�O`�$ઃ�k��� R-�قU�yS�
���<��U�CR|s�	���m��a���R�����dO��4�<h���X++��¤`�1���.M�ȡ��K+��������+��a�CH�|0z���y�s��\��=�~w�fG���4���a��1�Y*_�V[d��_ƽ�N� �Z�k���Zrԏ�f����|��uQ���m�}:U�q��g�|nm�=��y܃ͭ
A���5 PeL���8w+�u��h���o��4��[�����P[<�ۛ�����r��dM��'��'��F�8@�>@�5�E_�"0�g�$�n"�Ƨ�¸��ڂ�d@|��+�|�#<*{����:9mu��0�����Hy˺M��-��Y�w�̷�f:=�<JL��J�i�,�fݳ53�q#�,���_��|q�>���o�߳B�P�/u;f]WcQ5�i����>����%�mϲ� �S���4|���XS�4nȋ��*&���[&oL7�������5V�5����X�=!����<�Staƺ���K0hN� �-��I�+������כl:m@y�UX�q<���u�-V�[74�6f�,����+���͖� ~�&nȬZ��f!7�%u�A �jų�1'��.��=�f+�M�g��y>�'��걩\�?�������B�S[N9�V�4y�y���#
L�1cE�.煵P�L4�_7Ֆ���Ŗ,�a��T�.�V�M��k(�X�O�N}Z��8u
�On��Pi(�vH�	�u�k�[m�h��(*��-���
	�˕#�����X�����y�8�#0���BМ�����	?�/�	4Y���Jc�����׹��s�-v;��V�^GT60��/@��&�L-d�9:c�����M�����w��N hQq��U�NW�=�%�Ң���������ߪ&�i<��[P���q�E��Wy��U�1+
P3���~W�u�^�!pY]�K`��9v����^���b
�wT_�Ex�h��:��cjsu�Y}�O�{�Zwն�F��M�w��C��͏�?�j�boӵ}8t�Z{-���&E�!>�_z\c���K��f�x%����\�6����.3�&�c'��ҟz�N�k�[�[X�;pP�Kb���[4�H�g��LH��}�y�K��m�nn�����;���Dަ=T�A��h�>{���z]��2L�!Q��p���=V:��gГ%XOG��f�VN��H�{x���O   m�i;>�L%����m�;����C�V�"�������x�*�k���?5Q��;�t�=vc�C� �0�἞��?i���.z����k�q�.�b԰�c���y���a�UvZr��ER �NkO��R�sf�|�������b����2���QEk�gFc�g+s?'���<�^${�
w<�x��}t�Oza��R6͋�h�S��V1���J�c��:٢R�3)�-�&5N�qKݨc?�_�ګMt�L�[� �M����+�`z=
�id��l=�j\]"�)�v>�s�ұ�_����.���լ��R��`��M���r.�8�y|H�8�lg�`&7�� �N�x5��q_�>��x��?��ݻ��n�Ŏ����ܨ<���j5B r_����^���Ǡ��0[�gQ�};X�\��� �k7o(�|�^Ui����{t�"7��i�t�=F���,F� ����N��/���h�>�As4�<����׀╍�VH�-�eC`)�����3&�\�&�[���_�M��5�,����2����/�\վU�5�����b$�ȃezcR�m���7����|&�����1����+kn�~~���:�2��k�]0x.���f�ǿ�_�it�3H�@����IU�B���6�֒�<�ΐ�$Y������{����g�?f��[8��p�2y�&-޴���1	 ��A�v���`�9�t$[�^}�����A����#�6���>�����r��Z�(v�a�~�l'y����z
Y�79��|S��᳎�+�Ρ�Dqo� ���v�h����'� �M�O�jÂ�y'�#��fh4�כ��t�cG&�[d��s�~kW��RBQ`���߉��ǖ�݊���5	Tҩ����nɤ���8! ׳�Ԟ�{-���8r%k9��ߨ`@�В���lK쪑�A�Z3۽�3���H��>Ĩ8�`���9��PV?
�/N  wH� �(E��Fx�� �x >R����0C��6k���V�tM�R��h��|@�2�"ktNR��c����^���T�UPȋ�ߜ�����pِ��Q$�YQ�~�i/.�O?�I�.1�aX_ ���-h�<m5�?9=����{55eNCW��3+߀}nO�6��V�*$�c�I�џ^����v��6��P
���7
 ޔ�k2}b�?ٕ;�yYKg��a�ل���M���ZEU+6YY�"0����x {�?��<��9{	��^~J�jM"�9��9L�2�C%�X����-m�y��b4�5td���$9�ede���7`b̳Nɿ��u� ���,��ࡃ�z��u�~ ���~���L�B�t`����7ZwR�.Ez��.r/5	�2�������;���X�j��UxLt�6� ������+Ֆ&��X(��ja0��ᤲ�H��4-q|~����:e���܆�xg"ȫ�H�pp��և_w�{RYk�����P� 3ؚ��++;;9�\g����/�[���l��h/[.����F�Ȅ�0�7Ҵ�gۿf�6�Yv=��oh�K���k�.���IAː��O�($�S��tK�= 䖫�.��[|s�j$GNQг���?vo��l�xv���&�̑���`Uy:�V��[V�Bb��(/3�v��'���d3���EǇkU]��������N��2�|�u��0L}�Fq��:�8[��P������'��?����Nq�N�)��^\b��+5BH��`B�G�4۫ȳ��\�74�|T*�Cm�m&��2����P�GE���mfN^�q	C����i���+*W�7E�,P��3��_:��q��t˽�ҟ���kß���M��Sظ��ZR�f�IF�f�eD1�15,�9�%��ދ9-AڷX�A= X��*�t�_��;�F����)Xy�j�_/�&
\�FN�6��L���U�A[��f�ulT�K�ʌn�j���n3�]���*�����\�ZGh�f��01�\���[����S�cC��������w��w�v]�C���/�K�|�2Ӯ{ۿl}���/�m����T�F�KV�ѫWp��+��QL���g{Z�bhm�g�F_��h��s`-��D����pnQ�5!H�v�4�%z��轗�uF'�R�$:������{QGf�Ѿ��~��_�����k�u���{��c]Y��V�Ǒ�z�)��Ou'J�aC��3���楡���8ub�e��u����R𯝳�N^-���� �����(�V7@��\�Ap�Tm��5����-����H��$.W.P���ؙݨ�H#r<�#��� ;����䧫#aZyH�8�q�<3���2ljE�Od�.�:����J0�2d�J��}<���٤�̯;���Y�K�������hK��r�e����N��1("W엎)��N�Ae��А��
KF?�k��)h��-ƛd.�q��֍�_��r^�mg7��d��D���Ua0f'X�!�U�e�S&�z7�T�[P._zŝ.+w��X1`�U&��p)����`���E����Z��^�i�-n��RrU�iP�Ϡ�%!�����oM��L1�w�w��*/����O8g�	8iqP_��p��rHs�[9��2�s�n�^^B�ٶ�> @����9����#fb����>�[U�s�i$v��F�tO'�a7 ��4xp�b��J�r>p�.�QM��B��HJ�.�H'd�[���V�g�q(Vf[�]v���1��zUk�Z.[K��s�����QsY���
��f/��j ��������1�N\�U7�3�uz�����l��7�mj�ݹ���C�y���u�6��yo8�Dϱ�v��մ�D3��|/	�^�\�/�}M��ھXS�'����a�P�&l�h47lԏ�u/�i��탰20h�k�{����]3���>
{��!~&4�E:�v��ܾ�R��A�|��ln��a��,q����d��&��Mwl�2�7s���~�6�r(�U��m
j;**�~_3�t'�[�u�t����VH���:!z�,,��	��w��M�Qa����/)�%b�F�V�	����w�F���@Ė�;����	�����+������&H��7�U6��v���T�h9�� ����iu�(���XR�;�Gb���ڎ����Mk�o�0�I�}�M�E��㙥\A�I��8\�>��*�4 Y1m$��;[?ȇ{*)�K�������N���\���%`��	��%�R���Ȳ��x��`K�U��e�"�L�W�-T�q@ ��fY��+O�܁�/����L*��	\SKФ�8��0����8 P���Bd}���\�~��5di�˯w��fyx�t�1>"uioh�Xwܤ�Q�Ƽ�����\��7+��ۮ6��,�s����	׵����I��*
�4P5�܀���߄�&�?X<�7Xg���@��o_�w��Ch;��%
��`w�K���wi�-�g?s��j�h���y�|�x� 4��K�9nbd�?�N����D���Q|�R�R�͹1�]
1��wF$�����mf��#�,�	����~���^�9���ȌO=���Kx�l��_z���Yj�d���CD�4��?�hoX�5��	K�fa�2Ӊ��_�Q�����?s��������8x��a���%�eK	IS4> �F�J�����%��+�$ �ʇ7E���}U��\S�;䤛��B���t�R�!�ґzo�}oA��>՜Ev���lt���Һ�T�"�M�
�%ťP-�����f^|	�Y|8�q3��d�ɾT�oB"*Y�ky.؍����&�9�/A�<�q����»�gkg�F<��I��3��oa��������R�F�	�˟��X�1��x�q�����E^��Wp���V�3��K\v��5D��l�o�"�;Yz�
�⌹K�5	�mM��$S����qՎg��.z^~��^E�����F-��R]T�k���M�'�cH���Hq[pA� ��6+A�vd����7b�S"dϖ�p�M�#Ѐ�uq�#���J{���,S+x���?�@�p���9�Q���k��وlE�*�|�J��l��oj�4^R���G���׸�����1���Xmb�V�j ���헁VSͬ&�E���&�],f�z�C�S��;�������
{,;�΂��@���}=�0��刻���yD���"��W��@Ny���T��o{�tǟm���꒞R�۹� '�e0��2L��c�YZ���Q�}��4#�G<g�,E��[$�O46Q��K���J%{����;Q�� ӿ���g����TA���y���u���^>�W<s��b#ө���~���s}��X�z��(��r����_�BOx�J�f�d��H酦�=b�R�YS�2�A��E����/��_!�8>T�]}����-(H��R��_����'"eL.�qeWKr��?D�E����ȸ����l�q��V�=��֑���Y
���Ƴ��Nbߙ�j�bC��%�Ij@�S�>nRor M�E� ��j��N��Lp�Ѱ::Ic��C6�n�-G
w�H���ʠK��w����p@I:��\�]�J�����3�=O��.ԯk���=�b�=ŧT���Z_�vtd��kal��������gf�N�U��6k���fiP �JN�D�7|��hD��*�C�麍IDl�P�ϐ�n"A}(k�����9�'���t'7��B�qq
���[vt:PW녘e��,��?�M;�����iIRP��#�>�S�2����S�x��.����u�i�J8	7RL-�xOm�ZsU�wm��,�N^���E��/����&�vU�{����7X����2��f9�M���
�o=�� ��_�l�f�\�]c��<���-K|�3��`of�U0㓔�2����	=ܶ�:Ԉ�6�Yx�G-��LG0O��4�r`{��t�7I�=a��djb$}B<3Hy��I���nT���`�%����/\�o;9r��m]\��>�3�½�w�;�P�%���-��dŝ�������''ֆOE��m�5PK"�8ߧo�d�dΏ3�Ɔ�q�O�]��+C���j��ö!s��O����f%�ڤ�Z�`7� dE�g����$���Fns��;����4��W�N���.����Ʀ��t��RTO�VY\�,*S"|k۴���f(ЯN�b��w{���9�2M�7� l�T�6͵Œ���_��p�$���H�#nuD���J��{صzQ���B�jh�$0a�a��vTXw�H!o�P�F%���$���5F�e���G��<�pF֭8�}����1Px�K�PR�b��`���Wڵw�������t�H�l�a%��	���U6+~d�+��AT�v�[�����U
��?gZAyÂ�4���t�%�7�p�d�x�}��PPPH{���#Uj���vx����wx>p��j��*��z�h���U
}Tz�7Kd����ZV0�����l}��܇��Us��7��3�GŸ��aU��wxj�:���Z�!����$r��@0�Kv��|����@mT���}��:/���J]���d��Ѯ>>/B���K�.u�r�R)���M����øM�.LI"(�v�5	��Z �vg>��_�j.w�$�3t�Tv6S���W�&f�9��6Gɝy1v<�x�<:��(�֭�25cd�7w�"�7�`� 7��j�%��7����I�Q���Lj9)��*4�?%��Ky�|�Dlt��Nz����h!w-|0݌�	=0E�T�?�
�˩옫�MlO&�%}V�<f pG?���(�1ː�e�bӮ6��*�O���AN��]H���9O���i�-LO��=խ�nľ�����M��+ς�����:�z��n^������0&��������߹��\�. 1���K#ټ�������lA��<��T.?B0s�qa�&z-̓� *$Tv��%;K�oI��.�'N=wxj8�1���=�_8�&!�>+��ɛՖ���%��T�6y�%  ?
���n����9
l``���˕(cg3.!BAb���Ybܒ�<���;��28����k���v�TX#��%���t �l�1��h��gq��Sal���� F���NAAQl.��t��h.n��S?��4����.6����SG'�I���w�t�32ig<�{6��z)�:�(�YT姪�NJ>�e��c���C�V�9�}x7�㖀d�m��-~R��TS������.�y$�m��|�Op47v,e�b!������u��9��W�仲�ovl�5��wkG��x��ɷd�L+�1�m�:c~F-�$?=�Ǽ~;�,�v�����V�=�j�v"�"�;��cx�����׎�0��ܓy�����'˖�y��9�N��n�@����=R�Z��اx���vZ6'�%)�t}z�@f�~Jq�-�G�������`T[���D��z�"�`ݡ���sMƶVKci~v3�S=+C����h��i/c�-)�3ɣ{lWZ�9���$����-����UR�!��ܜ>'8�V'���̩)��4G��W�����F�5�d������=����[fIj#�n���|ǿ�R�\�l��X�E��6�ɜW�=��=	<?�Z����)j%~�"V���˲h�%�k~��[�ͥ�ڼ��@�ר��2?�s�+�+�&��Cz�N�~�I�I������#�j�h�����<2I���F��D󙤸X�Q��Fnدn�B����=�uY���Z6r�3z���6nu��exe@�0��BL}��5�A5Y�o�YEɉ�:�P���Y���$>�[tW���`O�t����e�h� �UJ��˵�G��b]V��Z��-��M�����Ĥk\���Oٮo?��N#!��e?*l+�:�k��Oy��ߤz�\�x�<-tZ�$&G�K?V��	�X>��^_ۡt9����L��8��J��  ]�	�N��;Q�R�'O�W�.+_��4���� @Ȓ�A:'f�t_{�F�h����YLR�uEc��cԹݦJތ��<�����{A�@�UD*�C������hȓ�0ሮ���J�6��D�̅�$Ng������S��'[�+���]�f�/*,����N�{;No�oB &��j��ы�y�O��<�*���m��`ڊ�{ݴ�אK�ˍ*�>�V�~q:1%w��4�l�}o|r��LIA���M�&���=,���C���-u�w��`�f����η�L��k����P���2r ��:'d���mb�R���<+����A����S`���jc6Z�`_�c���M�KF�u?��8��痋����x��q�yqF9����Vg9������`z����k��P|�/���W$o\��\��\�4�pP���i��a�I���]jn��>gɕ�#��ӎ�ി�[H���ׅ�*Q�]�����������ΐ�6?�u�wi;��1ݬ��2G�A:��\�t��Ē���]�K�>1[�4SPZi�_)�O<m�ˌ�_ l-��"4�F#�U��$�g�3ɥ���򲕃��V�Z
4�1`&��	)�t��ղ�@���ŋl?E�8�I@Ⱦ�ьR�7�]Z��D��Kqٷ�d�y q́F7��͊����;�4�ēӤZ�n�r>�:�p^�p�BQe����Ӂl�Li��w��H[���zW˾,4=,��ປ�6�0rE�+�12'�H�x��;��Y?�6��I���lX���-��!$�\$C��:@3/3�'+�����s��n��7]u]Wy�|'Z��\x��m�T%��VXI�ˀ_��.y�8*wjPZG+���?��]�!�s 5�g���so�f;4 6��RYUcy7��:4(`n�n�NS�߭6�]}�YE��'�s�����xMr~S�IO�9-;��P F�2�ks��U��>靸9���"?SOf`WY�W�U�W��C� ��66�����g�O��a��������V]��G��$ �H��5�Ie
�5�d��/��|t~��զ��ܯ�w��=˞F�w�1�秫����{�0�՗�}#b����q�	�[��t�����[��Y����ʴ	�������,5�Z�G�*0G��j�o	,�`C^
�6�`\�H���c�8{��ԫ�\-��o��ZKS̩e���Xe��g�]#)\�g}�	�R�������q���:��]&8�����X�A����o�� 	���j5䝩Y:�������#����+PihÕ^�?+�=Ae27�v�d�{j����gY�Gfx�)�R�"��P��,'P��F�[Й��j�Dx��$_��v���J!_ ��]�mG@��f�~`O���φ�J������%�!�k� �8鷅��L�㩈��ޮOYf���Kک��~����됴��qЋ�'h[��������r������_���U�A~?�<i3�h���x/��ti��LiZ�]�*�,~� ��mRؖ���\��L�V�
̺�~pV:~������g� :(#�'�so�T���ZK�s3�g_b����}�A�p�@�ƚ�^x�!緼��]ݗ��N8��P2qo���
R����ˇs'��6[��#��WΡ	���F��� W<�q����faƐ��v��l^a���N�i�/���oe���
JNw��� n�4�o�V�J��v§D<���Rs��q�A�N��"ʾ�ڛ�����UC��72���v^���_��_��V!���6m.�xN=�N�l��e���T�l2g=wv����G���7���?��3��rӌ�)������1H~h�����{���k����R��Z�~�OR ��:�.�kܭ�s�r�Жx�W���*�����[+aۊ�|������3mcxY>t��cO����h��z���@�(7�d+	z��Ȱ�N�$I��j��d������웈Q5YgC�Z|	_����:h�q����8��Z�qX��~y��f����[�k%l���S����d�@s	�9f��rL�?�n��A,�9�i���ݼ�D�	��� ����9Ɔ��;[�$�-�����?�k��ӑKLs���k$������%���8"V����d�JꀖҊ��zo�3g�ܙѵ��*�B4�����LjF�k����H5�A �󩍈4ٚ7�� 0-�&�p���MC��Xa�C�t	�Ʋ�����4��� 3jz��ٓg2s��0O�g���C�Ko�$K��:�Z؄�h��eQ'�����['Z�S;k�B��Ap�~�1�L�i�2PtSpp;�h�]��v�Cpk�]���Ƈ~���o4�Č#�4�����Z��� ��E-�wW�]�v`�DY�C"��+�z��z�������5�¿�h�U02���4D���Nem��.�2GI�w���W�>��m>
�c��<�ӄZ��|kS~�/Z�NA6�12�_d�Gű�q�\_��m;�b�m����6~a���)ǰ�_/6Ag�Wz����\�/S+<�xy�����*I�`���w���h��0V����Vz��"��<ro�,�s9F?�W�D����NgN�EJy�Gk�D�hh���`�93��)V&�Ƌ�̘�/.�LV����&�6|kVl�y�7Uv�N��C����*�J,-���w�G�˱6M@�ky�|�r�TF���ʃ�)��j:C������YM�$����N�O� /��1{P�^R�����0�:@6�c������Q���1	 �l�Ij����!�o�aV��Gobs�]������'t�?Șn�$+.*L�$���e(��r�۔z�X�J��#�IL�ېw+�g���c�t���3-�|�Z�W��i�t>PƏ�}�7����{H��*o�?�!�夠��6f����� \�E���ʵ���ȿ�O�# ���	�-v7Ť�M�i��6(���zZyJlPj@�pZn넬?:k���D�>�j�2IQ�1W$���KJ�Z�%ĸn�������l�.��A�/���+�rA�	�����=)�K���1�cLy��k�:X w�^�G-�p�ֱ�^�P�԰��w��1�����S����o�<>��j�&���/�i����8��)Eb�̷��wg|�/燣bN�g�1y��WARC>Y�r�^Me����519\�h�v�g��E������HM�Í�n@�2�����bn������Ā��d�bc}1X+�P��!��+ �s7A_m/����o�DH��Nm8ѹT��j��4����G�t��D4s�Q����� L;���I�W���I(��a�?�S)Fx�Y���� �Cu���HC��)�&��%1s_��(�����O��'p�/�����4K?1�#���B�P��������b �Io��p�����W���GU���Ǒ��� �{"<8fX����F	��(��##�+n�L��� ~�a��p,����d����n�����
k��ƒ��]K�P_�^}��{��sS��.[�O۟:�T3�<ٱ!�q�g�Vi��z�1�F=��s0��ؽ����g��e�OU��bs�<0�䶊�ItF��=?�@���J�}�;��5H������#��C=ܭ^� Mލ��Q��l/:p܍���7x.˔|�b%��q�����u�#��Y��$%� ��ϥ݁ ��/@��	�����쇁\�H6����b��E�HZ������3��b��..�a?1��-k�%��?Ho��n��eLW�b�Ƞ�6����Oo����Z��V(��Z���A6�<�8]�0�7�SCM���7g?=�,}�>�ǎ�)0�����Q�!m>m���T/��@}<�:�4c��99��>��b��}����}k�"r	lc5u�+}Cp�7 <"�^�=�R�r+ؔ��Bn�O*Ef��HmIm{�6���l��z�"�o���ns��@��N���
b�!�!P_�T����l�IbM�~T�3��c�m�]y1ce(>I��wS;�|��+����E����ƦW}2Qx0���!��O`V������{�j�R��I,Kx �x���nAe��V�#�'	 �k
o ʭ9���VE`�<T�6�v���4R=qU��"�iz��T�@�Ǣ0���/<e.�D�Y��)b�������qQ���ƍB�=�auF$O�4�,��O�D�� ��Mc�4��P��4d��&ٔ2m��\_#���Z�����ְ� ǇW��ڎ���q�:����h�L�J>[?��:
"���,f�Z�*���R�L��C����㦕{T�iq�N:_�acX�l�J��r�a�|s�q݉
-��i`�7o}���X�ԯ���"�.Χ����H}��ؑ"�H@G�n�ަao~$׋B�'���v"��eJ�-P�n��QL�և@���+%B-���BF~�>!d��p'�}��\�ΏKvΓ�n�q�-��h�4��>�!�E�����|`��ʫ�t���S�*������dզ/�x��,O��������� ���b]xL��w%��Jb�(�DƤqvl�7�:S��՚ٻYĠ>G�Gs~R7�w�@���J$�eV� ��وT��.]C�O�ł�-od�w��
ގ�|:�����Xn����:]Hy�I"��a�dZ���ڏ�����^��޹J~�1��
���*/9&�X^�;⚬����7��dO%�I���I�K��⍝m �V��A����4I�Fd�Ӡ�B�j���hպ��0œ2ح�2���.)L/��������ok�&��ݙg�p�d�`�L�2��<����Nw��Y��5�}�5%����$�+�2����#I�:��n�c���Kq��G{g���B�A�b6~ Mrrr�Y}���A��N���J2����y�݆���Ⱦ䉕t���v��񞫡9�(q�[0{:�޹=*�]��R[������������dٕp�87o��3�EK�	�w�4O6�����a�{�^k���N��x|o�E��vpp;cF!W�8+�˦ڱ��˫u2�S�DY�畈^L���_�Đ;�՛� �������I$�Gu SRLS�P�9���o����1����v�)s�+��<)��L������#q�%�=en�c�J���Ǒ�GQ�<�-O���B􇆔��/����xnsk����9:�Ḡ'Y�<=���mxj�k���K=��5Y~�ے�\���ٻ��ׅ�є\eb�i���2�i�:~Q�{~����38L8~��w3}�+$��� �(��+Z�
���s�*���Wu\�_'O���`J1�f?l��fX�S`m�=�[�ߎY�Mɶ�/I'_�P��M�v���F�G �枏轡x�A<���a���S�Z�DQ �'�4���8�>���.���:VVq����Qj�ղ��ٜj��I���`k
=���=���Sw�M�r�a�M�q���^�\YD�{��g���a?�>����&��H��D�}��R�zR����#0���%c��zd��c���*
X�x(Q�=Y� v��O��c_������񚰡sJ�aB%9 �迭�2(%�&D�"�3\��������ǌ�����}��D��Y���4G�)�x ��WH��"��j��kBZ����NS��5�˿�е�����Aܥc�778����6G��ŀ��nLL,:V��;��D�u��i�8��i��>�0���|�;0�F,�h�<��RG��T8]6���ԭ�ö́��C"�zC�V�o������$���Tٱ���
ƁNo���]����\_[��ድ�rF&����U��%�?^!�-Xz���i'�:8?���;s��(�ǅ����!��d�O���&d�7K�F}����6-9�7�ؤv>5M�Læ�J���P���Z�`������_�Ai'�|� "_������w����}E6����<���Rƶ�5|}� ���u��q�ʛ�7_&6����K�xiռ+���zt�����xe_:�,�����`����F����\��x
�����������ó��3� ���'Q�M}��3Atwu�[�#Q
��LD��Mt^li�$��xD�@&p������g��&"�M�R������Z�6&�� ×����^O��&��j)�=�o��0U�}o�mQ���̜*q���E��0붨r��;��=��I���$c�x����S��g$����7Á#J�׬�G��
�8ؐ��V#u�'@`U��5���O.��4�H	B@�����>ce���^��#sTbD)	HYf�L��]d��,] '��-������Z�U���Y�o��������9N@i�kI�!IL��w�Bޛ*�E�w�.d�~�}�g<J.v���!�>]���1�;��qb��f������������5⟙$�2'�����iʸ!���u��\��{����^j�S���%��DĈj��R��I��F��h��1��������\��{�	��;5inM�����| �d�����j_�'� Wt]���ʰ���-����AP3�4�����_6�T2����Q�ٌ:|57��͍�z3s[c�n.���,\�˕DN�����IT|D��=q�p�{.���(���i��Kk�ש(ɗȶmW�g����g�v&�0/�^AMq%H��:������nf;�̓/�Kr_��W�6m�_1傐�XK�%2�t,�[LK=S�-�=K ���aN��T�����Z���F��c7�C�-�K�:t���P���?nt׿}G],��}�ӬE�3R`6�dd�������İ	�n�2�O��tc��R�8+m���2�-��{����>�wq�[� 8��\�`Ĺc.�
�3���'`��T����Z������3�0�E�p�孰�?�x�/�����z.�vhg/��,���\~�Ã�l��ȥ4�
g"3ʏ�(�������8�U�F�H�Y�����ru	�(nv��LHm	�x��5���D��(2�h���]i$���u�s?_'���O8*q�"�ծ�G�1��}�Os`-�t{ǃ��6l���ٸuK|�b�s�ސ9E����B��(&[b��ǂ���̓�#�����#�<^�d\��J���H o7�-�t��'�z����Py��M4�k�-@��<�#�t���G>I�7n�?=]���(8��[���aڔ��= 8X������{Ud��_�<2��iH���MD���gxc�Q$)��^%0pH���ȧ��F��u{�c�y[r�1�_qtx�4ٿ�\`h&8�u,X�06�~fvRU'q����v@�>��j;(̆�K��N�wLU��I.���y�6fw)�Q���4|�_��Ĥ_�U_�AT��R^�[]�&Vji��Ӵ��㠋V���_��U�0|�J�?�t�_�Sxby��n>��1��� Լ}H0��RWn�JY��U3 a�uv���L�̒����?���:��	-�Q�gh�콶��9�����@	#��9���x�K/叏���@#̂x�87g"� ��?���|����G�=��g����k5qm3�}���бu^��(E�ɕ6������{��I�K�nq�&/q��!���>��՘�0l$��R3R4٨��uߦ}�'>z�@� ��xfD/�Z����;l�Ům��'�,��g��|��Z���(((���"�����.Z.֒oʆ�uq�B��Yp�����\?_��_���7�T��T�a�%/�h�K�	��pV����;��x�U>��kC��"���Eӳ�ߣ_766�o9L���UT���K���xJ>3�>و��\�A�7�l�|��J�6�ɬJ���-޲K�	Ln�%�
�^B�4L�����x�z�;�]n���D�ԁ�{}T)���(�|C�>�Y-��/��ڭ��j("���S�jؘ���fW��e�N��G��*�]A�i>f����\�e��ج�1<mok*���i$8��l��Й����Td���37.��\�+�:����\_���.��ÂX�hI!L�&c�%�
/_���)� _u'B�L��T�"G�1�����%^��A��;r��}�gn�ߟ
x������=[�b�:�b�W��>t�9�fݞ�|t�BB9�VVj9'vR�F�m��:LǋS��y�U�d�բ'�l����7=��f/����omz��g�CfKي-��P�HN��#?��)�Ai<��!?� ��\D:���G�z��	�sݦ5
�QPR��e ���ـ^�� �H�42����*��GlQ3��2��I|<2�Lh�(���y�����RgLQj�2��PO���3LX$����]�[M�J�ج?�A?社Љ�U�"U��V�����[�N߉ğ�n��CK>�Ũ=��y��R�6�,��<��o{_�h]�ܽ���)�#R����������|�NO:�i�4�V�o��6���-VL�O����?~s U�2�)UT6�A��۠�޼�UQݛ�N�[\�3r�1Q[���?�Wjg[�WnRy���q��Go~'�bX�D�we}Z��o$��FE������4���>P�f����u�[��$�O�>{����x�攀?=�{@�{!�J�I���N�S<.W�N���7bz�R�7�6^�E���i�cQ�4Y?��&e4��	jub�N��F�f�u�("�^1f���½�#�T�|�p���}�=�e����FC"�+(<�p��;�~��m\K���ǋ����N�b*�=[��
�u�M�w��L@+b���ຳs�j�h��/D
�GO�쾵�6(ST�UU+k�0	�����k^�Ɲ��6��pd��+�Zu�(��*�*�������L�5�9��/�5y��֘bI�o��ru.{s�f�o��>���y�D��p�s�gsZ��@���9<FUϖ�V=f3�R�}���Ɔ�ir�*���ךSQ�NV�o�~_;ݶ@�v�����Eă�\I9θ�I
��o
�e/�hh)��V��U�p��Dù'�?����<^�{�$c��xPY��1�~Lm�N�#�A��?O�-��]i�.�v�M>r�x?5�t����\XU}}�O�Y��5��9j�'���fG��� (�;�z�1g��ZG^H\��5����짟C`[�o��v��ѡ��Ce�����J���Y�Z���3���[~/��4(�7/L�IFH]s|�H\;��Aȃ����$�/�o�d	[�T=���:���JȦ�jX�*e�nCt�"69-�g�V܏u]zY�?����:Kt%�3�ɽ��H���q�/L>����+�����Ͼ��s�ݭŕ1M5�ʐ)3g��/B���`��K��R}���wX�@rl���[�=�$b����������rP�RR�������c6��a�Zb��-h�]D���p��i&\>�Y�@$w&L�l�gp5��ݯG���[��K2��X�<"��.r����
���(!tV��-�ϳ���j!�9�Qv�`M�-����8B[O��!Y�M��c2����fœ�湥�Aӌ	L�+�T��M6�gR� ��x��G����Lض�ܥE��ab��a|ɚ;1C=�wY�O�]yX�� ~k������� Ws[��=n�o���&�����|~�9�ԡ�.C�'��k`3��[� m5��m�w���[�[P�%���:�ͧ�k���N]�٩j�Q0�ȁ��sEXр��(���z�O	F��'ݫ]��`�U]��I�զ��� ��+��&��q�(Y8~	���W����2=,���'2�����������~oa?�����G��¹g�:;uM{��]�^��~����\ �:���'x�((|х8^�Awd�o����*�~�@]N��ܸC*4�X�_�%�/�O�\]'O"y��S&ZG�x��$�X�:���9�WL��S(܋�� ��ڧ���x�����XB��`ÜF8}8ĝ�T$�'��L��u����9
�P�r�U�����"ְߙ���Y�}���;��޳�uՋ������N�~"�O_dG��͕��W䅉�n�vŘ#����#?l-�5��H��+N�d�3e�������+��T`j�~�u�c`]j���9�G��h�Bֺs��Ȇ�ܡ$�>2dvZ��$�å�U)��(7��z6G��{q%��7S���4�{v�����i)�Z�D��T�M�E)G	l���X����M����ʲ-7Փ+�wX���sG��5�:IVR�^�dHG_��/{�Is{t�O�&�k�=��d�f�SkQZ*kk���5�w$�Be<�lV�m��P�i{��LٟM,�zLS�,���xu����F��C��P�{��l'c{�	B$�f9�$/��%1ӇBEV\��b����^i��1/F�6	AS�~7qF��Y�vz@��~����dt&o�VzP�,��=�
����7�w���+���X�� mUJ��7Q�'2����ǆ�*��> 
rBgD
U��[���4��ߞ�����^%4��5�d\<���<a�u{����)q��O-p=h�S���2`>�au���e�������z��+Hn\.�s�_�Ș���A5]�,�~�$�����W'�[�2�t�':�R1ٴ�<��{!��D���ڼ`Um��<xDo������<i��-�lZ'@^�T%�Rܧq��Τ
D�Q)VH�P�c<�������� ,�a��d�K2��/(���2����������-�,t�������k�%6o3O�8[o�\��)�`��UL��,F��B�ʳ����s/�Ҧ80�8ŷ�Y��Mh���g7l~�}M L�,�>�:*�g#$�|U>^�*!7��O�P����P;����U~���򩷊�{����)�?ePpIg"�'w�^/�~4�<1�a�<}��r�*~D5���m���g7�.:s9ɣwe��GY-[�ٻq����Pw���q������Xp,��n����l�� �^��\D�����⅒>ŷ�3����I�쓶���:V��t�c�����c6q�U��T���w�UF	��S�3yL��d�@��k�	.Q~.B�o�����A����CM6!���̕Sq=7�����㋔�X��-�a37S�Ĉ�����>w_��o��KF�5~D�Ov���R������	딑;���/%��J��gk�-T/Чz��-<Yʇ`��B����;&���呤R��"�
���sE_�������nC�C��et��is�� ��E9	�ps�{�%�6�Ht܎V1� �޹�W�5���������=�PQ�ծ1�����QK���0�S�O�J:<.��0O�;F�&s[�j8[芄_{Ƿ��PL��w
)𡇂|�%u����~J����g>����~X��
�G�*hY�F� h�H#:DܞI}��Qe�j~M������N�.E�f��-���]�id?�ǩ�ڊ"�z���
�S���<�_�c��5��@�����\��Gu����.ۣ�w9f�-.y�QCv��M#N?������̣�gR'>ʺZ|����>�2�7Df!���`�%ُ&}�.���ڇ'W����@�_�W޼Y]�	�P���ɾ_?�H.]�=�!����C���W��,
I���nn]��,���_�~o��q���Lw���wu2ўbea��V�[
�#��wR��T�\L(�a��/�����Hj HM��u���F�婾��cz�h�{�iYƝ�_O�&�M��Jn�f�:�����+
�Eq�Ɲ��� ��	��www������A��Ki��n�#��s���>k�U�jι�j��?G����i��[h�R��ԃ,��Y�������v�`����-1� �ԭW9-�\il7�Qj��e[�~Z�aX5=lS�n�mQ���;E���cH����'[�qw� xv��.��g��/����N�kV�R��4\��4��e4��l"�|+߭�F���%�+/���H1�[p2��U��k�j	8;]eA�~mڼH���bR��E�2�}̳��߼,N���&��YA;�:5����^����~��>ܰ�d���h�^�Y�OL{��1��R�~��0��@}Z��?p�/p���R�}֍�g�җ��P�7*��(�T�����C������:K&���$�}'�g��ij��T'Z�Քv�Ci�.X��\So*aF�;�Z[��0���k�Β��D�]�N8�<z�i�T�]��&����$�/�����e4������D��m�H�|���0��"�ԿVU�Ω��w���6��,��yY��zeЈ�E)?�3w`ӗ�V�c��֟���r�Z�t��^����Z���ډW�S2�O��{1Q	
g:��ܱұMk�E�s�F���L�xk�m�ԫV���
�jlը.���YK |�OU���� ���SA��Q�$�7ߊ��7%����`+�m���#�2H!���o�BZ���aPL����J�ٴ�:��8��l���6�/�uT��f�a���;�G ��N��=X��.@{���I�Ci�TT��?nptuƨ��2bP�38]޽��8:pi���F��u��7@�I"�������ܙ��ab @(�����P�s���5g�|� �vCd0�iP9�9t��~���FJ~\b��l��`�/ķ�O$`�iE����5
��s�p��MՆK���6�'^l;o�
s�ڶ��s�RJ���G+_��?�m���/�#
��D�\�L�a��C���	�!*_n4K��DTn��[M�]��)G_���{���ut�����S\0�#���Y��=�8�iJ���N*ͽn������Ql��*e��P��h�.��_��2���OU�����e�*ƣ�Uč�F���7�R�=�g,+7�O�P!E��O��s�~�v����T�PP��k�֦����-�����(��M�<}���OO�5�N����*��׎݅�k���| &�����%%j����8��c�]�b��?v����,��^[�a^ܥ#��Y���ÿ��#���w&��oD�|\���=�������ļ�ï��*ǿ��D�$?��t��~x�^���.�h�5^wʶ�y�ƟE���T_���s�U�3�W$�!����v/캤��d�l SN�6����/�:�
��ցߔ��Ĭ���k��g��S-:N��_XD�HDk�O�f�<��6�����n�n|�4�n��+XI�aT:X���6�M4
I3��qk?=���#TA?�RM}u@��O��Kc��eO � +��f�<g����l���4r)l
Od�}<�Zo�Q��������eÂ��hlZ�����q$ ؾq�÷j�WɊ��zVy�L�kSd�@ɠ|��C��~��hq����_`�/}��O]��M�/=a�f��JKǩ�+�1ų��F=n`� =�čf�����$ͪ�'J�'�Ь����AIN��"�Q�pk~���MfI�>hի�X*�S�6B6n���ښ�摺ʕe��+�kȪ>��p`�
�������T��U�i�FG����3�̆��|Q�P�UF��(���^�3�5~4�Ɉ�ߺ�5��$J��GK"-�F�&��L�}niUa�3,�op�j=�pݸ%'2�22�g���9.��A�a��͇"ꤿ��at��E3s���ds
�tm�|-{Lt8�-o�f� {��4�1
�`������.��hd�A���?�������E��]]�X#A
je�A��ONĩ����V��~,*svk_����9[�U�:OWe�!�$�{�H}��ָ��At����O(�RA��?<�ps����h��]�8��j
�<q52e�qZ���'��4��K��|�a^���m����F%lh�:~���1�<�Ũ��N��[����ԁ�Cl`v�XP�sl�~(�u$-(��aT1U��1������Mԥ�5͠�oA�_g_�/��N�ޔW�K+�0��Ƿ��l��k�Qn�D�m��u�f�|��:,����$�6t���0��NH�a̸������I^�4����c��������_;R R:n&�@��T167�j�e_ɗ�^�
.���{�<�UU@�DJ��'B����j\5����I�k^a�.M#�@bҬ����̬�X�L-�q�o�:�9�Y����k��s�6�@U\��
�;�n�l�q����R�|cڪp^U�f
6���⒖9�G��T��$�i�敔������Ƅg���Co�eB�d׸�7��{��Q��F.%��f�$����[A���w���I�������[��k�n���{��nӒ���|�Fq�
�� �����H��LH�i	o-�G�z�mPkr0خ���$�җ��E�1�?������4+h�kY��6��T.�|��O2Y��L��*�c���jP:oPw������Li�G�<r��4Ջ�e�VO�R��P;!!��W�Ua�9O���t��v�o4��&\��Fm��|}ص{Lo��+�֯� cHWL!��Pq����0�/p��q*���m���2���Ex�r���YV��P-}7���P��0�T	ɻ�9mVh�����M����"���>��/劆���3�=}�O�����
��v	n��xHn���~/��{�D����~�hY��,
1k�X��]NW��x�� ܧ�mVY���;&[���w��jok����� �Q�Q�����r��T�r��x��@�Eѣ�d����s���ǰ^�]M4_�"�}�5��S���Md(�e�H��w��Ğ�Oi�\%�U��u�)���ǻ6���Ѝ���#�������I�3���z����%����(76�K������"z��c�,�J�[bG��ڄI�L�Gk!�V�ZO�߉�U)L�q�j	�k�w��G��Q�`F�t3�}Z$�#QȞ�,L�.�*��T�O�o$�q���$�7N�h����j;% t�",2N�Sm��uH%�	YV����o-{�=Cޯqe���}��T��Q��P��>����*��ƚ%3JώF�E��I�j��[m�E�lwİB�\K���WdY���H�T�<���BG�������L�J����l�ܖHL��&HC����);Nh*��P̤'��(�Yj�`2���m)M(�xF[{�d�nQ��^+�M2[�?��v������"j	�n]�Č��������<Oi�01�:a&	f%�U�@S��%�����تֈ���z�=,1����f΅L���=�P��u3��f#��TA���N��"X<�D�I[��C�(��pyk��;�i��\r�!NS9{|^4�AX}""�����y�{zM�˱��C�)��K�21|�V���T�EZ(:X	�<m����U�bG�/`��j�C�<�L��@�:��l�=]���Ho��{wse�t9$�I�_r����Ũ	J3��s����wp��-�ȡ���4�� I_�|
p�����)��u��~q����HVeW�XZ zڠ��N
���D�,�\$���'�@���Şy���,���O\�n�����`�iy��7�eX��竗�,�*�D�~hʚ�3d��qwF͘a�������!\WGJ1˚�͙g1[c0��۴#��ův��6.V?��e� g�<�W�����v��ZlJ3U�6c,��N�u����#�G���4��!]���`t���\�"�o�v��-i:�R� "1�����\��Ϊ����]fqB?����%)8Wo��mߠD�����sc�e�y��,����`�z��!���.�lQR۰�qo�X�:����Qi���0֘kD"|���0�3gi��1Aa�T�Եt�F�3�O�s,�n,��W��_�����P\�ы g��%�hi�M`ȹ�ܴ4���R��k����.)����wO�I������xn��_����O_���de?�mX��֝ۧQn˵�(���Ր�x����4��B4E�<أ���'x䄶��Ӣ(o�ȷA�r����v���ٝ����.O͈���58
��|�2y^�2��a���������x���w@���Lϐ��+=�<�ԭ�XK/�V�w��/e�u�L�k2bj�9]���9݌�\dm�5s >���T��ʔ�Y��g\�D�~���:E��e5���S�껿8M�ό������*��J"���\�^�+�M�K	q+��M�Lb!�c�t{�ҽ\ߒ�,D-��Jx��}F���A��s�Ѷ���`o?����%���"��5��<����x��Q�mɮ�*G~yeը�3	A�W�����������P�k�G1�2�.�,*�V_<��^D�K��ySN/���Q�[ڧ�D��!\�����PG��+�I�ٗ�)7��}\�/��[��Ǹ����*g��d�}����k���.�}����tuC#t�)w�.覊�N�r���w���f�V�	^c�0&��SQ�/{�
�!�̨�p����{F[,ly�o�������	�\Ÿ�\HBbR������w��R��ǳ�#@dI�R�� a��z�Y�jnk%�y�-�`A�G��-;�iA/��k�A�M(���R����P��1�M��/r�vQsj��% �O{n�������*R�-�a�֦���`�L��S}*K[�JS�)��Oi�!�}��>�2Kz�߼�z��p�c�i�h����wq��=�/�,e�	~ttɏk:�x��POط/2�3t�BD��Լc 8�v��Z������$d*�'���ЩJz�Q�����rx���whm	ye��Ԗ[�LC	a��ew��nR�?8���CI_�.R�M����!xp(:K&4�%�^+`�u��|,L�}qL���9�R.��5~�®f�o2��@��*a�:���%@�`"��(��U&�c����wC���Ć�2�5�@���yb��}��lޯJI ҉�*͉��$>�&�B��_��T�c�k�A2>�o�׀��O/�Y���ڥC�ȥ_U\k��^O�5����jd}pސ��DkA�ӻ�YB��F�k�7r����*E�l�7kp�8����e�����-;�Ǵ��;�2WA:��fT/�5�]>
�ǩ)���u���Z�	�`���� 2�����9���ϻ$4O��6�?j�:	_�k��?�O��� ���n�ۉ����Ga$�оj��`�mF-3,��B+��}�Nq@�ّ�{Xg#37��z������hr��k}��� #�hW�Q��g�s��v2 ��ĵ<Ez���ӓ�-���ae��m�|��i���YN��;��)��Kް/�z&�T���i�z��4���������g�`)1�Cs\�1��fs�B�����Ʀ��J�Ӵ@)/�-B�����U��|MSZB{����/�0�&[D���X%HT/�eu�x�&�f���R���˕uj!�	>^#��u�� �A���Q�"~ס"�L�����)t�7\^��ܫF��HTu���b鄠�GR�7Q�~��:[�O�&�g�͇��"i�љ���\�[ai���I�C���P|O�OZ>F��vV!Z݀�*-%[3C�:�;���yƿ�^���)��ɀ��~q���S
A����:�f��~�W�4�\��̥�̎/��G�J�}%�*RB'.C��˞M�y���K���}�x�)
Nj�J�,y���������N/���Zz�S�:qW��D�2(Kմm,I��H�5�*�կ0����¹1HwlK�h#�z��p=ō(*a���2x��$g��.Lĵ������̃�j�|�蹓���7ؑ����|Aܨ�M;!����R�z����?!m.�ryO͢�q��q҃r���+K�a�p����(�;�Ȍ#�OcY�5��Z�_�b�	Mxp�jO4��Z��1���&r|s���D�+rG^&[�>5t~�qѸ�XQt���v���	x�i����7�����u}$*,��=��>!�~���?��̭eY��d٧��~Ϲ�pKYd'�SSz�y�y�h�,��9��&�;9���'MB|�ru����|s���z�b5�e��[����`Hӆ>��<N�-�M8-v����k�X�s�c��_lǪrV�������dòJY��'mF�<�����]%�y��g � K���t��ǭt
�9� O/�k�"+M��e���
13�	��O�xu�աl��"��%�[8v���RZ�6���ϜŁ���b	g�kN>��t�!tP�z#MPBA~{�̤炩�}Ef���f���t��D��4�)�T�H<&*���vK��$�K<�]	�"K�=��o̶�w�/%,֠o�O5�o�t=���N�LK�V&2y�o�<��	&6�����eϳ7�C�����ʭ,�2�9�ߤ���|�ǹ6-Sۦ0�g�8��!CKL�K������v8�O*+-:u�"wcf.��H�桺��OWI�Z�O����l��'�9�N�(\�g�Ƴ_<$l$�m�HK��0��y�@�Ng���9eG�swy�RoW*edrR7Н���{�w����U2�$�������N�H�T��� �בsZ��-��o��k��_׳�&ӗ�U�=�Y(���N��@�C0��Q�=˒��U��<]�}]�t��p�r�D�d<������C�ʭ�0h';��s�t>W�Ϋg��ҵ�>��~2����w�E��E����ɕ�-����!_�|�y����Æ����э��`ߟ���Af��V�eP�h�2��S�Q�\�wo53�]���m��t�`�������3��2u��ฤ-�\u 2�Κ'S��9��ԇ�5IG/�],qR�}����@��Ӽ\b5�2�Į��o��`t�tx9������3��TI�n����B>4YjF�W����yҫ�������ӽ�;�
rv[P�p<gx3R�"����[��
cKV�\<�*�:��"�E��[�} �pn|W�c���3g�bQ2Z�f������+$�&d�0#��A*�{5wTm�&���-��`��3?,��N�kӣN4���)��$t���7r���Ɂ��D�g�B�1߳C��_N�2ok�n�ٺ��ɑ�Ky�݌����'Dծ�a��9[#�5��s,erP�������'#V����w�[Ȏ�*�h�Vz+��A`�4����[�������[Y��	��	�3��������v�	�31���^iR�鎳qv��Ev�Bޱ�ćW:)�us�e��D�"���)񭀿���x�ঢ়?��`��%��j��kEg��k�4ʒ����i�y�Aw�t�������%owcN�u�9񛎵����H��`t���yS�S4W��q��h��fu7ΐ#O�?P��3�pn� ⌯2��Z�%_����'�<���������������UOq��K�d�}�߸h;#�8yٿ��_���ȟ�؇�\3(�H&���kS�������l�����^��YInk�����"0���P���[��90i�p�El�pĂ1o�r*m�H��*��Ciw&~�$y��/U�{��ͪV�O`a����B����=Q��@7�pv�(Y�4��铳7JD-�e�����aðI�P@YB�&��� w�we2ډ�r�|��D�����E]B�ꏩ�6|-Yl�.c�Dh���J@����"����˦Z��Ӱ�nu s��A/@���l��𔶻���i#aЋ�-��37�A����OCӅ^|��h�s�{FJ��\p�-��m�9K-&\��f�A�\O{]�������s���5�d��O&���i�m2_��˙������z�F���ǋ_x�� �ʉX�-�~��5����\9'����F�:�����	y6?����j�`�Qrz��O�6�Ap���"�v�5��>J�qc6u	�9`�UId��C�g�ީ�]O3Hu�-'��O��~a�ǯ�@��m:~'�b�a`��ّs����}��c-B6�� :q�Y�˛��]r=a�Y� � N=q�І�k
�����'�"��<5��X	��;V�K,qv�HGk��S���a�$��'���/K���X���&���[(�6ێ0������=@����D�ɱ�}���[�۶�qMɧc�G�8�f����O^3Ǆ�x�m`BG�0�٭�=����@��3[�To�ח�dv}�>9_�V�a..�7���<��Eۀ��)��̫�҄�$���n����W2��10�Vva�ϣ���3U�(1(�T��;_b����BP�I�j�� ��
�0�ʦ¥�2L(�����n�]LĈ�,p#�B{E�c4�j�%kW�_-��*h��{��^�|���,�2�����Ѯ4}!��'m@�^?>�����>�gv��ٯ�)-��ւk�Y~בa7���b�0�p��U/
3���i��;���1��g�v�oR}�^.r<�x�Jh�ǱO�tL�6VW-�$cP�{-���������ߔНX�0�g�;�LaĒ?ov���M�4���s����z�����4z�čZ�Uq�=�)$8t��ц�>�G0�H�^ҹ�a�m�jt۠��u��ڌ*k�������hjC Ls���W)�xW�_!�z����fI�'�����|��jq���RA�=��U��A~vMg]�&+p[���?8����h�M��m@�	��Z�%��ecBYp΁è�'}������F�����Q<���ZB,��5۫�I�S�����n("�C�}%���|Իd�3o�Y��jT0��Iu��F��L���1j����Q�}>���_�#�E�%���^�5Ū7���߳�(@r�O8����L>�����li ��*��ݨuz�:��64X�+P~��V:ۈ�/���1�	���kϙ���{��$��:,H;��k�a��O�1�{���+�u%bXvm�{�; =�ɮӘ�7i��r�7�߭h������xh�5¨�ǫ��>�ҁA�&D��Ih:�����x�"`9İ�h��5fzK�ܬ���!��yv0ꑹ����33��;#ճ�z���1�7�V�K����-���J�F�6t�sl�%A��}��+�I)�s[��O�꭭��ٮ�-7�{�A��9ש��?F��x�p���&��RZz��(p�%=	�d_7.E>	4��!J������ǒ74`h�e$i�2u�kѕ��/���n�A)�&#kD+_c�/n���v)�,����[��nN�i�s�jJ����a���	�c��#����Od���i�O�G�dƐo���&X�˔�fx��p�w_��N;�zĊ�|M�y��Q��W����E�x��{YI���/�~ڄ* � ��k�Ǝ��R�W���tj��jA��.�T���(m��ə� �F1������QX���Fy����M�ą<p��>�u��:�4����*fE�
�&&F���j�qR��qzE
q����8���7�jy�?�*� ��k-#a����{o�Ǹ�͌�Z�A��"/aT��|+�:Fue,ٍ! *�σc��L��*G�ĦϷ�?DL�.o���h�N`9�z.�P�ٽ�Y�n�����f���w��:� K�0��2DX���qm�71����9N�X�!o���r�=�|�]C@���PX��㐔�E���$�RǍ����~����Ʊ�r�CK�ظ/�T;b����]'r�qa�(��7�(	�����@8U�|���k�֊��[���}��ؗ�?�M#�n����o����7�$A�"i/{�������6���.�G�'�6b^Ƶ����!��m��j����_��K��;��������Z�h��sq��P{r"����v�_���/�@��{����n7x\�9`��ʞ/j�ct}���~r56&��/����Ō��uQ�7�����j$̼=z�֍s7~�&aP��	 ��hj�kQm�I}�|� ��ʲJ����	�)HL���3G��#�6�S��i
�j�t�ymFcĂ'$y�2������l���X���/�@���ۯ� x�4Z��ʫ��6����0�tߐ��K�W8�3��k�y&�;u'Ǟ�)��{:?�V�{-�~@���,x����֭��h��6���HC��?�e���x��I���E������>u�̌yM��<�$a��y=�]K^ K]<1q[J%�R�PzX���c�ݝ���W��g���od��Hˇ,�����rgH|��(:_�� ����}g�L\<r����4U»=m��,vG~^K���"�����^�_�����~8�?�N�=��%�/���gh��nGa���5߬��k=��Dg�l�"��I�=	����38b��$��X�����4���
��^Ж"T5_*T&�!��c��Q�$C��B�V������[�z%�y*/�.5�J����b�UblHQ�My�Q�I����m���(�i����}�c�3�R?��]�h�(�"5��J>��(ڎ[�ˡB��|ڒ磫.���~$m�
�y1;��x7J .�>:?���5-�7L4�ey+�5�L���0ʘ����2]���}��.�F-�MQ�	V����`��|���p�4î�� ��z.j��$@����!nuC�|��������`[��SPa���V��2
(n�#����XB�F�Z����9��K�7�������u�@.mŧ��[O�g�a;��6����������5���@M�ٺ�,8V�ưJ��ro�sDk����I�\lL����g��Z�Х�PiۋI��.n�,��:�l<��&�"�ޠ�1����p9��ğٍ�(��0���bYY~7^-:ir��k�+�I����~�_��O�NvGq���,�@��b~�A�,��MM&FP|�� �85J�,����gF�p1K{@��6Q�VI֊���n9��Sg���֣ԋ����	l���р�������}��C�8;�3��Ǐa��Jy=]��ARb��A�=��_hd�
�t����*M����\�5��g�#\�0DZ*��,�nғ�}%Q�vpO���㓬�=ä����,`��Q�ۇ E���r�2�m�P��3-�F�Nu&��w_��|����D?�CI�n����
K��P���q�I��j�Q�~%0�p"�~�P���h�]��~���[�o�\眼�N=�Ġ /��I)�Z�,!
��0sII)J��'\3&h��T��wqJ�Co_�d�Ҩhg��`� �2+���d��m�*�M(��D���=lb�3;�"_9A��S&t%z��!:�Q�v�(�2�9פ�*wal�"'�3L0q�a��+��S��@��aձ"�1�I�R���^�Aǜ8r�5W'ag�E��i:o�D~���.�ri��(_�:�c��{�4�]��od+�[r�l�Zz�o�e�M������m�4��������va��̢�m-��Y�ܛS�32��T�D��{�%RKZ�>67��4��}kD)��f<����$�d�����l,�:=�
�\˿�8\&}�hU��%-��PV�x���0�:�`��g?�l�<�+p��0��u���ɵ����w�Pȗ����� ��������&��娰췇�y����"!�us�����:�@#0����%�Vvl�0?�F4��g_���@3�y�k��$K�DW5��7c�Ғ��]��ǘ�v�MF�:R!�u2E��,n�y�g��L��� ��8Ħ�f&W5��.�ڪ��6A�]uv�p}�z�rQ����HG��)k�~�.�F��m��7C�\��	(�*s�ð琹�����D�0�Ez�0��!y
��.��R���_���96X_F�ػ��'�c����<��?J��<�����^�LH��X��ΰ8�62��i�4r��Hx�_Sq�V̋���fC�Х�����KB��\�m�_U����čZ��Һt�ek��,ݶ �G`����5�_҂�����k�T�③�!:�_X�φ�"-��#�M�k+�ԏGxg55Ȏ�A(*/�#\�$�#���E����O���������Q"��������R�� ��|%UN0�4$v�j|��7���S��b��m�Q��
��,b|�`�+���s$�D�% �2�{�8�T��r�R��ᎫV;����0��&0sg-x�r���or�Eœ�]���Q�A�{.sY�p�C:rWb���?B��3�s��kM��9��k��RA��Z��iU�5d-�E0A���|: A��P;��8x�e�\���{���C4�GU&7C������L���ꏗ�����H�k7^}z� `2_˽K�]�����*��b��.�3��Q3���.$3 �ف~I
Z8�C˘�\�9�+ʁ��8̻R
i����d�X;�n��8�/�e�g�H�'�͓a�WA����l*�օ���ےF�?v~��}y�id�%�V��&�Z�����Qx�����Q,_K�s<��9X�U����	8w�#v;�7d�h�@e��g����)�� w����̅1�I��@ԜY���/=�[�s�.�2�Cnf��:��U1��I�cR��3z�"{��������I�q��1�=��:����eA�j������p�nm��{�BC�J�-��-���r&�պ�mdҶ;���d�We}p^�ǫ�"�=��V"O��'̮�u&����S9�o�9_������Nz7�wzl��
X��TJ�#�O����Џ��yԌj�]w�)�R����xq�F�}�t�[G�`O�?wJ�����"��������LMc�5�@��e���+�����."�85�T��*����;�0*8K�����|z�������N��\��E%A��7mϱ���q�gr�[�ߝ�n2�8p�~;Y�fN�>:�=�d\#����}���%h�N����#��|�nѬ3��$�|1$3�oka�ٻE�i���V�
�U�_%��U)}��<�����ek�Tkb2����q_�O�.�'�);����mn�N�X���A�3F�"rL��6�����h��5��4���[թ\OQ=�V��)�h��5̯h�T�m +Z��hg�yRL�nz �����C�����y�<�	��������c�@�fqK�[�n1U��!�(V��q�h��E�]�1pԿ�EL�7��be�D����I�}�^rݑVK/��3���j-��"��L��G��<�����NS�e�(Q1����Q#GB��ҥQI��N�B���x��?X�[i*�o�	��ŢK��;����`_Lh|&?�C���Sk���)��~�>��s7R �rx���F)�\U�������և�d��vG' B��}��n����D����)_��_H���K?��ۄ�O/�T��\B!P���@P�%Sȳ)��bk�&<�ճ�!Sb�����h5�(�;�5+��΀$QS�v��2���R��y7��(d��{I�{]0����|��?DӾ�Ι���m2����_7*y��ut:ǘـ3e)W�_� �p��WM���5���L��RqtLB���+žJ���&��5�%�:�t)�����%�3$�
L<��S�<=5�yh���k;�����$��԰U�z<��G�)dѴnkK'#?z �ǝ��S��^����A��	�&i��K3����ý�P����2��ǵ"�$���jt�@·�.�Q]j<=�|���*��	�kEhq`�~��]��nd�?�o���5��5x�%ĸ�~M�d
Z�;������'�B�`�Zn��(/����j�7���!s����:Qt����2��h�Ox�\���Ez���`��u��4��3�$d�%~����;���MAR�E�T����Q��A�x�׹P&lN�MU{�K�p̨�ga��P�]h�b�̯�9�h�<�C�VX�(�C^Yg�=�8"�|b�p��X�|�����-���}����7'юʊ�?Cȱ#R6���o��.k��!(��!�tl$��uL\�ѽIVܼA#���%�*4�DJ�M'�u�Y��h��x'��u�_m7�-�@����T%�|��s�y�3O0��1�1O�%eQ�<�8��<q�6�/��bn�~��僻@�ᗱ",b=���Y��le�ޠzB�R|w�㑫W�0GZ��m�h��շ�S���Z�H��/\��0���v���`ٕ&J�g9l�3��p��� hp�Ю}[�59�����������s޹*�^�Ť���;c�3�@=KC[?���W�f䘕x��3`�h��wա�,0�y$���[�ξT*�z��pqڶ!,�|��Ar���t��]kI���Y���å�(����/�2㤥���NK��e��A�����[�ٶ938�����%��q2������C"�OJ�02w.�~�1H�o~9�|��\� ��E�XD�3�z�?�S(l�J�U�Op���h��$��J�ִC!$�b��^Kcc2���M�723vL�n��sp!?I�La���J�S�8w��L��������&����|���@�kG�S���CTG}�cr��9E+;�4������-�"o�=�~2��������t�D�~洏A�^�!�[�
��]���T��9:��]��dm?@�a�����Lc��+��μ|�yｍn�6�.�h,�>���Z�[o���R�a��gQK�E�AM�-�<.��GV\+j�#���Yo�C�۶�#��_ޡ�3H$O�&�TE��.#�~T�������?�>��R�P�2M����u��wȭhC�@$�	�5�������i8����d���/w�e��G\N�"�Щ<iJ$���n \M�[��d�� C.Ο�E+�יd	R�о�]O��x��:���/��١�5�(;�'p�)Iq�p�!��'8�5iq����񣕈<�.�o�ڋ0Ў$�7>e�VK�đ�鋭��T��~-�>��T
�t�����Q��~6EBٛ@ӃU&I8|��5��e
D+S�!������O	�����irN��꫇鋚��X=s4S��rz�z�iR��^���Y:��j�e��b��0��k���a��,g�IJ��&Gՠ̀Ӂ:�����z��CCm�C. 7:�lC�s��PW7�K��4~�G���t�<���}���Kλ��x�O��3�1���n����o�,�b[�QBɺ���n�{�RAx0���3��c F��틤g�5'��׬w�M8|yl�Q��-�.�^)��<�9���Oܲ;�N/����lʺ��Adu�޸���
A��N?fl�q�O��do-�	d�W'�4�HYd>"�-Οك����0n�Y�~�e$V��p�wX/)ӄe�Dr�ےX
�[�e#$2�Sg��a��/3g�^j ^>>Ϡ��N��1oe������^Sp��W�Zl�~�5/�)=SO���.�>��c�$���R�X���P��+�> ^3?���1�ȴ"5����y`�HwoP��	Xd�nn��!1(�
ZI���
� ��|g�sHO�A��O�J�({�=�p�;���4(�*j�����u��_�*����Be�X����ִ@�*�tf���_R�OB��Q�+Ѵ��
s�셪sP�%&
Ӹ�^X�!�rM�@�K_r�������,��t����Tb��U���p����O����7�)݁`��R8����:�t�V���'J:�A֌�{��'i��Q_��")*1�۱�7�-��m�ֺ~,�?�bМ؛�T�j�)5�9+�׮�"��d��Q�CKy�+�S��v9w�~����i�}iN�w+����a$f�#Aɀ28d-�M���t��ےV<߯w?^PN�,�k��7	E�4x�j�X3d�t�'~�i�R��H���z��d� t���*�#�[����ː���21˭܈��M����)�XHd�Hk�b����\�7��u�����us�Q�Xr��=aT.���ugi.�6&J��<A�R�7]>a��.6��O�	hp� ��������-�r��ڽC������-qA��W�(�S���+�V)2��t�*g~b��5*$��O_�d�����2���	��ep����������ܝl�����ڽO�p�����>����
�����L�%��� Ү���w�:�q-�eަ`W�rJ��C��j9/���f�r���C��`f*��Zt��ߔ�l:a�a5��&�(����^/�A�Dg��<�>�����
%��~���إ�H���[{jhQ�'h^㰺�>�C{��_�zC�	��Uz�x"����qOW����9"�la-;�X��-��?��AgۼL�)ɈҜ�������s�0���l�H�
@���+�c^��� �3M�B����a���ZI˽>BȒE����������h��ԑ�B���0�����W�[��p��BO��]�9��g����I	��K�~�R>�mZ᯵o�?e&�ѫ��1����`w���y�[���tP�PW����q̋���2-���tx��5��9���.' �Um6w����
�{�pv���֖��'�8���:��	i�=\=���`�:I�V�0��wH��}ͯ�7=��������un0 �2��r�~�a՞�Uj#���������c+��<������ 0i5M�а����A�~ǰ[$���X\3�ee�O(΋d��hݭE�ǩN�[I9�n�����U.c�χ�ͣ��v��1V�v�� ��1.|�>?vg@�� �����!�]��e�LM�
�< E�B>�'x�ȡp����r�l���R���qxj��f�6v�(�:���^�_�Y�[A�P�HZ�u$`80�G�Z���
Pu� ���:�����sD45� �z"���a<��Y8���.o�;r+�@PFl�x��t��s���*�����}��c����L�G���E���/3�la���\T�a���V��d��sT()(���Ǻ�Z���a:���G�(�L��@�B��z�N;i��^ ����KwAy�HRw�&j�l��hI�!�� }\���t�y���>j��I���8ܬҐ�,�c������{v�� ޒ�ȧ�,�p�^1��ٰ0���;�h��T�D��JѶ��\
N���/���y]+H~.�1X��x˕�U&l4���L�\�;�T�	$��,Em�Q��jtI���o��9VAAX��Wğ�d�[u]����P���(zQg�k�����^� K�0;��eϏ����n�����4d/��,��L���N@�&fPz�]��5�;L.�]���F�@�G,���k�O��0?s��b�YcS��]�U.k|���*{:�J;]��ن��Al���Q��^��� ^���9��\
������ٷ+�����%�%�����7f����<��m��uz���ou���a��F|��\K-ݑT��_g���%�2��ϫ�qz��k8#;�̸`o�A�~���o�tB�Xd�g��x�t��jqMO֕�l��+{�����/��i��(J+j��^��J�e�,<�:���^���ZPVd��`,��~~h�(��>#_/k��fT���;*
6�c��4g_8�y/�m���}6�f�[�t�-�=C�<�\�;����r��N�����fc?���r(�i��I�qhJ����M�H/�&�g�5߶[�ӊ=�3���3���3d\;�4���2��B5Zd/8뒵@�c02iR�-֧�!߇�b��m�M��="{ 䇳G��p�Jy|�UJ7�o7OoT�r�x�G�O�||b�2�D��~�8��I*�gd�����W`j^�w��M�[���+�!���j�N���?G�
-�`��=�;ZBr����M~_��4����c��eԼUꀊ��_���-��P��aMZ7��AC� ��
�W��0^�0�vd.��� 圴�k��^�~a=ܧ���q�7f[}���7lrJ�/D�%,Q��g�,��O~]}m/p�����LU���#�~\��$�wæ� !�HHB���a�y0i�ʛht�
$��.���4�E��{f�;Mi@�:c'���'�]�1�������(l�R�H)s��# �=3�{\�v�h85WF�N�������^D9DN��Lv_}�g���5�5[W[H
j�t��?�͗��`�0Èz�/���4�QWյ��;�O%�y�� �Y�(:Q�~LJ~��O�����	�X�M����۔�&4v��v:M�w�\-O���܁ښ��¡�^ࠨkۗ�����,0���L��R2��?k���`��P� ��f�M_Ow� g������(�^�|�Z��q�/��΅ց�9	���d�j}6�5��̲��� ]79��6SHS����[��U����Ɛ0H���賌B��/������[�\-�dB�+̭h�� �x5R��������G��Xр�Rϔ�_d.j��%�I����S�a����)��������
̢���+b�o�V���ʡW9z1K�)��g	�%�D4q�s���xe�j8�;�x@4�ʧ�b*20>��8G=��}����)L�݀�9j��~M�b��߭������Q�c'q@��p�\�*��'��^��	rk��T�� qE]w�7&��#�l�\P^��<��)�ً�.;���ǭIF[�Q��Y]��s���`���%"@ͦ��zy�����Yr`H���U��R��������RkOk뉣�C��'������ښ~��ẳb͊��ܞ��n�Ļ�� J.�IQ��&$�S�FI�~�&bWE]�9�MS4��k�ƍ2�]��(��@�y�P/���"��k@�,��B��U��ӎEZ~!�Ы	]� �ƭ�h���\���8o�������$��nI�[�$���M��}��ciڈ���]�M��2oۮ~���:��,� �� �q_#^Aqĕ
ɢ�K�5C�s��D<�aF�����P���1;-�og�p���\�*�N��KH��f�^:��5
�9�i�!Vҕ0k����ߝ-(�et`��{BE�iu��l1�R,��"���_�|3�]������l�]�BT�u��I��Wu�'����/iNIx�qaD#�z悸�"�Eth��(1�1G������d�}?U�l��;���}�(Uj�*n���iSB6�E�+�9�I�6[�R�1�Y.W���n�c{��(�yB/&�	�[عW���iε�h�)E+y�
���#[q��X1LQ8���@>YM��ܿi����C�V�{B8*�P��Џ�����(_f}�ї�[`zH����H';�*�4ْV�� ��Q����mW��`vyr?'�i8��*M�Q�8?�_XbqàZ�eZ��EW����*�?�&�����V=8$�a����)2Ζ��0��ln�[s�ѷ��~�*�Q���%��Ӵ����z����_q�U�Jz�%A���;S&n�n_�H�Eˎ�wz���9e�����7GI�H
��W�[���j4���{`�qn�����fN�l��Xmw��Tʨ_�L�ܭ��J�I3��AQ^���. OM]�W�4��r����0�t�m�e��,s�&[�k݉�{D��]n�ѳ���Ҳ�6�);��VZK�h�&�*̱����`����"B��|	�\���q�Ä�z	��Xʘ$#����Á����13���a��৊��(�@�����e���F���w7�*0Qq��?K>��3li�@D�aS��ѽK>��H8���m��4�F:��� �җ����E���P'u`LB+'N}�Qrq������A�G.YW3l?��~I�ꧡru+�����W�6�cJ6)�Xz��<A��/'�Y���m2�^�=�HZK2��Q�!Q��cs�q���k>��e�y�υE�+�Y^VJV�#dm��0a�)֚߿���^Ĳ��+�G�&����qhi�3}{����SÑ��ƍYayU�3����aR��[Y�m��s֥^��c��,J��8Ҵ�a,�/�ط��=����hZ������>�k���t�7�p��P�����vv �`�Ԝ��n�c�8_r��Ȃ�S�"}����~	}�!�c}�:mDG�C��Ɛ�?�-��	 �^3m�G�-z�Д��)2Gc�p̵j�m=:���j���2�l)fG!�tpbgm�������q�PI d��t2N�Z�zhcn܉��Y��GK"fj(���E�✐��A&�7����ue�%�h���ي2W��b��ΫM��p��i����ptrho�P^����0�g�-}�Ht.�D;I�^��
5Q�[
)�]>щ2�6��.2+���w��(�u�p���U�Z�}�̿�҃7pBy�pn@U�rl�����ҭ���~/�n��y�>��O�������ޯo����Go��q�bߩ�ze�ʌ�}_������1e#$XI�c��B���Q��m�0��Ȫo�|bR��0�^k#������(�
��PY���[)_���d)������X��g�ϑ�_d$��UNgQY�s�FR���'`qq{��*ф�˸�0��LiEZ��U���r���I�{ӳ�S�i��^)T�+K�un\�_v���7<��	��k>D뗐k�%�Ow	��i�S[�P��(��R�W�Zp��W?�L��vQ��o´���5�\ 0|�9	���<����� �j��ɐz�:��U�Ͳh�MN�|�Qf�ab���Rb��ȑ�r�%�p�4` �W�:���'À���J\�atE�So��is�EPw�At�vv��Z4H�-���Ԡ^�n�����x�}@����	eG�,�hE�1���|VBcZZ�X�|Al�V�y`�6=e����Td~������t�}e[�%��݅��P�w���mK%8#����g�J҂f��L")�h�L ��a¼���A�pD��I���ͷ���X�8�~~l�(�c�=P�V�Y#���½m��0_4^u��DP����2�����7��2	�����1E?3N���U������a 2�K
{2-����[�U��/=��A>�2QHDg&�4�Yko�j���%h�����(�"F-K��ўH�~^���)�(��	���ΰL�����f�e�%� �=C*<+���>��"�
4�|'��D��ў���8��	��F�e-���S��E��}9Qӝ*�h����I���=[�i�\�D���$��`��,�6����	�v(3���� 
�
#f#
��-Wn����B^)�kf�� �� ��A�����?��~�S��a���`��QH�25�Dl8��8��8iȧ9o'���}�i��΋N�C��u��hI�S�=�Zڞ֑2�B�y�bM�35m�)n�\�����7=�r�R��v =ph���r�oVz��i�lm�5�톆#@[��	�)���o� �%௄C3��AY.��&����׏�J����m^� ��{��:�{�5�M�{s���5����,+����;�$��ŀ�P����\��s�M��&6��j?v�l+·w-���AQ7�)�W��.ᚳ�n��n���1�D��	���Z����{���^\�����I�3t]'ƃJ�@��:w}y���Y�12���.��Y*�9+:,�PW*�P����a,/����w���N!N"�P�K��`���V�ibN��O���w�!�x�0Of]"��iy�죉�/9��g�]��j`����7�%��c�9�V U�������,��RͳF�KӶҨSŵ�ð�"�6g��RX5M��.�����֭��t E����5�+��z��k ��#�Qe�k����_F�F���[��}~������2/�ԏ*����A�[ӡ���ѻ��![MQ*��w/���B��1bO�4�TZ�dRF�$��T^o
�����N�]8�������O�^�f@�4�\�?�9v�a�ٛB����x��m�����@=]]]�йoa����aM�.Y��i�t�Ȱ�����Urr�u� �k�������ֺ��ʱy{��[/���=���_7�Z"Ş���������쟪T�����n��ɸ⑂l�Z�Mv�ޮ�W��#1�x�� �u�R�����aV�,hC��yG������4��ϳFD�䉫|�\4o�����p����J� ��#��`yB��-�O�(^��?�?��0���R�"��~A��e9Y[J����C�ݙ�n�7��#҈|�h�:�K��A���G���A�=�� �k�(�_4�^Mi6���+� ���0����E��Ȧ�ց�:�g�i9�~�ɤnk3�F�kG���v�����rSD�r�;O!8��v� �µ�����xQ(6�W�M,���'$�P:]ĶN^�;/�	�ԡ��v��7���A��$��+W�u�#^��œ��s���K��ë7C$؇Ed��
���?��i��T&��f$�A�L��s]������3�1?�hW�R�(4aY�*��1��ݢ��8���G�t��l��Ox�ӍIt���e� ;�Nv8���4��M��<I�DU�+Ǒ�'Cn�"�1�P�9�M�1Q�)F�3A�4D�	I�GD'�IO�yI�I�'��/��O�2��j�}�~]�=���6G/��ّ�#�Y�_��R��/��]���x��ȵ*]��/ǖ�'��Y�Ժ+ރu9i
�N�$���N�9�m�A����3���>�0ݡ�l[r|q D�|S��0[.m��)H�c�e�/�K�i[�O5�6�c�힏W]���I�%������gh��R._O{PKhK��k��*hן��� �\�c��l~l�T9��v��:��
c9Tg)�-P�w�<Gy�����n�ф�j��U+C��-�� \w�E1̐g���h����L�h����T{�IE���E!�0=�bQw�;�T�q���<ha��D��	����rh@w�]r��mPD��������Sɗh�Ȏ���G�bz��_1ոǪH�q�Μ����l���rU���E?�ZJw`�d���9��Ґx�M�� �غ��r�����"�e��d�<�F����6��e�4�܁|KC�J׹�)g�:,�����w{¿':;��vZ�[��M�~�N�n�7a�1�F-�u�����P��`���X�*_  \��h�&|������mW�K���m��c�G��Ҍ.�=M�Oe���|Dt�Y)��Y�?D,4ec����]���^A51E���Cx��xꃛ8�ȴr��X�lw����Z;�"�_�}�.?k3ʑ%'���z��Ō��#-��u�-+K
K/���O\[���Y�� �Xm��K$�bģ�����~K�$G�q#	T|_�j������S>�m�d	��a�k�3/����!�`�T�����}����B��p���:���l��� {D�v���W�XF�#��+�l]�Q���o���W}�N��M�"�U�~aw���m�8�C~�vT�����$���k)V�A���+V`��QRP��_W��k�.ik묪 �<��&�ø��]�M���9|K�{�zuH)���3�C�*`��0g��;C�%y%�@�Ւ��
�-(}g<���躋�Wd�Ei<ۃ��/܇���i��h ���T�X�������{���㋇kĬ���=�[ �*-e�v�4����Fu�i��<}Pso/�4�!������P�	�<���dz�QJ�Аb�	��VB=�%z(�2�=Gc�pN@t�(�hS0�{mR�W(f�d��|�*q�{��,���Q���n��L�c*s�6��	[ ��	�e�c  8���l���W�� �e;�N�t�Z�QM�������Β+ɠ�1����h���`����C�b���L�f!�t|ڪ�3�y���{H��z�ٿu�7�&���S��2��ԥ*�����)���"�w*�z�y�C(@m3�5M���\;�n��:�/#�1 �z�؉!߽���T�ۚ�����䞨�d��	��Q:|��yb5X=w
�K����'�[�bN�y�4?ƺ'�
]��=Y?H���	<w|��������b�F�yN`��a$D����q��c�?Bm�l�R�As��-�)�ol��̣Rn�����l5r�H��&��хc�9�L�9(.���%zFc���P�r�"�z�G� �v����D�;2!�N��F�� �X�|bieq6��̡��8�%������G:�dY�f§X�J��=��;!<ut�����u��":�j���^S>|���
�Vm�_̧��t����}���g����D�q!���60nsM�8��1��$Y>��BO��xi��|�Ghh�$w�h�5_ Q�y�R>�:�+�����]Mϊ�8;�-:�M�,(�?��]���ȄZ']�]qK�&�1Q$F�=��b �^֮mD���g��v��^3�_]��d�]�o��q]��M�ګ���RQ����xp�P�|�������fnMN.������+uQ���t�b���v_f��:7+��zH�<�e�(_b)�S{�چo�FS�Yl��	�k�'�7q������b�>S�>���~�=l	����T6����/�gT���J��w��.���Ρ^S�e�?�d֦=bry �}��+Ll�����#t\��.f���{��HOt����l�Z��v�:���<�pi.1��gY���o�)�P��C��d ���t}����i�t�7������a��r�,���V��1؆R���ԝ�5u�wc!g5,��z`M����oޫ@=4����+�e����,�J��yD����ʨu�K�C��h�g���h�~?����`:�5g#�`�쥒L�^vL�h��d���(�Y��uE��C�e�A_*�!���Sw$�C��nw`!�H�cMw��'#� ��e?ҝ��Q a��>�
�w�c�2�zVּ%���9VqnA:I���q��	:ِ_R��F��LK��c�Ў��t���<��<"?썆�,?ƙ�PWFsjPP� I�ۖ�i �yą7�Y t������(�1`~x+h��6�015��Y1�}�,�Eq��o�D7�{FJ�o����3��q�ޱ���X�b�%@�2`y�����,��O��Tf�U��{�-���+�!6�s�Ⱥ�b��&حI5��0�d�.h����_2�����qC=���0V�}�~r�<�Ҝj�lnF�>)��u��`���#8�?���9z���x�9O�a{Q���ѹK��[�o	ƒ��n4)alK�� ��ϐ+-�׎]S��/��h��X��r&��&�����e��JU��5|���Ԥ��_$��fy$�B���� |Z[�i��7⿚ �+��Қ��Xt^��ĥ�~M�T��J�P�$m��س�����=��\,/M���X#���(gc$e��K)�L��b=��<�e�0n�`.;�a������r�� ��6\b�9����2'Z#f��{b@
8&�# @@�y,R�+���/'��!�,f��3*O�s�<"47?�M*�C�.����ݐ���Y%�TmF��=G�9��K��!e��vd	�w�e�f�<7.��t��q?��l�G�k����\��>Q�!d0�������wk\-) �uR�P���oɸ��Ș�|ϲ�`��&u��ܷ��^4ڞϫ��ҙ	�
K�{�6����I#)���A�p!վ]�Ӌ�����io���]G�T_��sCEŖ֍�k�g�
�<��#!2}Fj�;Pi/�i�/uFH�>�ۥ�_�k�8�9��ԛ鯄���-f��0�e��A����џ������_u ~|�^��C��'�IJ��ׅ�n|�c��4E��uߘY���>�yH|������ I���2:i�M9�ܫ1"�*�P\��JH�@o�rAtчNzVR�+��.d_�;��S��X�5�/|Ńz�ހ��;�Lt��v��[��pD�L�r�d�k�c�I�^���!����^j*k�����[R���ڞ����oL%T5�-��z�C���4@�3)���l܈��G�T+i:F�����j�z�������r8��M��o��[�%�`��2M�(0�C��wseE+��;!8��G=�7��Q9y�)���\3x�6�ޞ�OF��2o�8�h+���'g�BݫVsRui��.Z͆�tn�'C��32�[�|�GPs\�rC玀W�)���*�@+*H�ruFX������l����I�M͕7B �#<��+1;p_�Y��+��˘��3ު��%�&Ю�o��(����km��X"N���X�in�}�����t��u�|Xg�u�2ka���u�[H�6�q�?�hD��LC�I�+4�����K4��A�4Y<:)��^;��f;�mV#4}��P��%ҮnI�O9ؓḑ���s�`�T���h��~�q}Ω���!iХT�-c~����[�$�o��9��6#@k��������	}�J9����<��KxY�)�D� ��Q�~��ng@]O�<�Ƅ-�L������9tɮ��o�6��1
�F;��6`O4������PK̡2S��g�n��G���ٓ���S��G%x����x��Ȉd��ߟ�3�m����h�ݔ�:e[[���~��(/�(�v ��Ð7ʭ<~�@i"]-N[#*��=��d\�U�)������{S�z#}�^��;�:?3Ԡ�,�^Ī��I�Ex�p�I��]lo\��N��˧��c��1&L篜�����^>N�0��R�K��)�^��d ig��i��N󴄜�ێ�b���+pw�T����X�?8�@0H��*����������,�X��$�����$���h�Њ��i����vG�0vtPCb�Α^�~����i"�9#$��i>c��3��/
��Y�>���Oi�q �x�]�0�%�*�[��uk������+���L4�<�4���CP�G��>L��=�Ӯo���g�JGq����D]�W�5�u�ކ�uJ,C�ySr�W)�>�1���A��9���v�m��v狭"�����L��S����?��J&R�e\�2uf����Y8;����}�j� gX��	��*��]&p�{���N!&Q� �ה�w>�k�}O�Ep_�r��I�6�vHa�җO�UF�S�-�N�%ۙ-Et"48����U߀��lk��/�V���?M��a[��Z&b��,��JZ�Wd�2�`=�6��X��M���vޓ_�����	?ȡ><�9�J��F� �#�~E'�M��l5��'�2�C�L�~������>� ;� w�f���^$�\��+�'�ۻ��D�l&m���O� ˚�Uیq ?#~�9��j@y{���FvÛz[z�/��
2�~�<��g3tgƐ�������Ө�\U�|�l��_�X�R3p��t��n�K�1U������_���F��z�gh�Hb�Y�/��D��8\C�.�
j�'���8�9��⒀�yO~jǘ�Y ��=HR:����
r�Z����9H��i�N��k����2�Я�ŷAX�y�x���k9���Qwҁ���+�[o�=O�6����8�NF��n䧥�Op��Z�UE�YJ�u�B%<j&��p���8���D�O�Y�=��'� �ٿ��Taڃx���&8�j�>/��r���n!������N���u��B�����qصE��	3�&���y�઴���య)�����%K)��DF���L�x���HJR#���sH�?h�t_���Ш�B�˜�,��I���,py�N�=�P�B��c��S 5��vS���O��|D�ǥ��@�o:��S��=�S��5����){��[n��c����)B�foe���u_e��ǯe9�e�T"&��?>�>ʶ����~���{��x�j�;@b�O+n�S���Rҽ.��	�v``��*��k[/��D8�,��4v�b/ ��)B�1O6d�ur��a3�d	m�(��U���/���jZ8���iP�����"?"�U;|����PaA����Ҹ*Rb%����@KB���}����/�o��H�J����*�[����跼4�*{Wx�zg��/n���Z��h8�e{�Ì���Da�h��	�����=�&H��u�9n����ǫdb����y0'?�4�?fS����sr�����C���-c��٫1q��o�!7�:��_�>���o-�_�^)4�	�`.n�l�0z�=���O]O�}Jی�&��*�T��Ǧ��}?��8bN���c#�|�LzĘ� �� ig��z�d��\�?����V�װ\�(0��4]uw�\PpG#f���/Օ�j	I��`)q�q�˗?Q;�����RR�Ƶ�jK��=�S�"s�4
�&L*)�-�rkh�����9��r��w(����s$�e@���^�X
Æ��fq�&n�o?��6�R��/��#yT���AC����p���c]q��/R���X���ѭ�=
?H:a8�H6��T����p�?d%���j<Z�����ۏ���lRC��x��̹_��W����p�Jݩ�,W���H�Ș%1��&��)#�T[�4{���T����)���5^� �V	k���zz��rA�{G���p[d�"ߏ䨅v]>�Ҡv���)\Ky��(Xmr(���9����0gB�[^��}|jH��E��#���V�!����)��,U�0w��Ԅ�^F���|�g۝	�䏗k�]Otp�%��8A���?�j��kHک��:F�Qi�z�H��9��}з��_p�
��o�(��"n�^��a�����|��%qBg����ף$��%J��Ӵb����|�G��	�����R-@t3ec3�{l��/�쀷���l�����(�U�-��T2&�|rE�m7����هr��_�Dp&��������n.Sҵ�r��&n���=�xS�ކE������b��I�qW����3M~?1g���{5�{xϢ�#��L�?X ��2?J�7N���i��z�J����)�Dk��"��-ܼ�\"-��{�Ĥ�p��}Q����W�O�����L�@�+~ԕ�|�1��[�IkL}DA֩ʔ)�\E����{|�F)F��k,p?�m�M���X�Z��2�D���gt6P�G���o�Ì�MJ�l�p˽�8��ߖE����k��L{�8�#A�����l�.�'��l��$�	�ӂj��(�?��^���Y���<Q�h�a{�N��cOS?�r�G�����n��4C�^l�T���겾�ʇPq2=�K�.������"YD�^dv���A(�F8�ׄ4����3����K|�CH���e�:�oɊ.����\*Ox��,���!�8��/�R�_V��K�U�~�h`����B�e�F#���b����R[{&�u���8k���2�a��� ���L�F���R�$��
���_ w��?�;��;���v�I#��^]�j����^���}�lد^b�1�6ҢR�X�^q᭓廧W6�S�I؋�l�;^C��Թ������al���z.�uѯa2o�13,L�sE5i�OOV�3�^ͪ?��f�̱p'h�U;����ed�?�����xG��{�'O�s�sJO��-�%;��@��ƺG�{A�ļ|bqv�}��R����s��!�h�f4u�A�\�egһ�X0��8Џ����ٕ��1��q�)r��ff4�!��Z���<�GRj�l�x�l� K�C�]h�+�H>e��yJ�z�,�f�c\�+�}"���s��?!g�w�Й4��4xA�/����5�[v�~�ՌI����I���X���8"�G�3.S�d]ݧW^|��A�1�"%����{hR8�=U�W�b��m�yM2�/�``Z\w�0�����t��i�PK   6f�X	�\  \  /   images/898ac7d1-13d0-4a1b-8b5c-ab7066f4327a.png�W�W��%����K`鮥;%����n��I�EV� !݋�t�>��;�̝{��qft�U𰩱  ���"��:��&�ߔ���'X^���  ���q1��w��S2���t���y�s�p��z����T�|M ��)���YfO�����~qv��ّ��v�C�m��� 91��3�,.���3��2м�P%sVOV����$�\09�U,��Ka�����fv�6{{l����c}uu�ڻ����\"�4����h�v�Y�!^����!7�)�Nʑ��[��������y�B�{rrr/[��q�$�|g�Q\P\�_��m����?���Z�|�}�X__�-��pM���������O{uNF����0M8�W-�Դ��۱�茀��4�7�/c���'ˎ�{ƀ������ka��r-�v����}|/}||4�y}>~�w�R1)d�-�uYvW��������kkkW�O��V.nn�� ��|'��I����K$A~���:���0/�j�ڍ>�^�,��ۛ���x��krΖ[�2��������I����}b�t�#���3jL�Tp�f���%�M��&g>���h����Ŝ#)}V�c}pr`�A�W�rm('���� � ���0���7, ZB��{����p_�u~�>55��ŗ�L7u��aMH����euU�򢻋�@q19n�ViFq�{$'��Q2��SGv�< ���Z3?d(9_�S���'���Jߧ�kc���h���dNF��1�;U{�K�����B�~�o��JL��S�d���b��*��+f`uy��[!s^���w����%]�sCã�~�����������x� �r�fr+�T�^����>uMֵ�컁1t���!��Y*��%p�fWD�����Auu�]��E�R999�e���R���M뭡��'�i�=N�#U�LԾ��<�ۯ���g~��d,x�>�-�&Inv]_���]����*V �|�������B��.{��,s5��D���#��Y�]��f�h,�2�@������?@=Y-���犸��{ǦvFϵ{�����eI��<�T�ۮ�?�=����#D@c]�!��Wg�>6���g�T��Tnƻ;� x��ú�(���F�����.Y����֞N�;=��U�v#�Q�EA��� ���o����T�����<�]Ц���P�U�X殎1��ٽ���ş��z��ɿ�eN�]�jGs���\{{�0W�5(���f��,4��S*��A� sIh��Nw2�J�l�ਜ਼��X�2h��3x��%Ǩ�j�L����	!Y�@�G�s��*�l���#�ie�	IM�f�� �����W��D�����<;a�+~"�
z��;B�t�U�ť�&֗ff�1ɭ�}q��2JZ����vj�6q�^ c�Ì�M���(�0E�⇥�<���-��~ �*�塈(-�?���Ć��$??���q�yr!Y��:�	�7�M��m��;e |F]Z0�u��Ӿj\pW()I�+)�F�8epr/a'?�޳����]_А��Y�5�����ff��Eig������G��i�	��7?���y���yVq�]�x����
��1�fs�(�/�s��l�R:-���^(��6?�s���N?���eu�-�&�i�czkH��Q]��"uj�Fz�0��a��5�f�H�EK���c/I{k`��pG��ߥ=n��[����ڥ.w�p�a�a*h4�Vb%F�J�觍��vgc����<n�����a��eG����U���A�5��֊	w)��~��+����i�f��uaΚ�¯��k����[ ��陙�.`ra�AlqC�h����6�S��'i���nSo�'�$���ٹ����WKF~�!��%�0d\��Em�O]䃍��+��qLi�\���k>
;|P��&�Q6P40L:G����J7>0�e+��f�Ԡ���,��{*�$��Q��$h��#��~�i��*	:�R=�0O�!�������d�!8�۠( 4����U��-�l*�L�� ����\���ch�*���bh�J؆*�m K�1��JM;���s��¢k=�{�5���l^6�&cW4|Y}}wl��j�i{�y������Q�S
�	�Jk����rl(@�%ݴ'm�ڕm~�����=�tLV��%0#)��{C��@Z3��h`��[�0$/x�t ��g�?�H�!�B�tV�+61��BG�nna�R���o�^2�J����+�Oic6|������$��,�8`��~K��	K������儃��{(������v�>�)�����'�ςE�\���udJ�HG����5�ؑ\J�M���M����D[���#y���� طt.����Z������C�+[�H�����nK!IG~\���@�#.f[��=�-�#�=	�k�T����B-�m�7��p�������'��9BL�[Xvل��Ԥ0��L�;,K��Rd�n��5���,�J2^�A�+*RR�����g���U�)��ݗU4�����s�c������Fۦ`e�m6vX�t����V��X7��������F�M���1��7?tK�z+~>�\�鑵z���.���il0Ͷ��z�����o�j���W�)���d6p�n��X�����5D���'�((���W�_��r�wu�5��b��ߏ�7{4����۔iA2�x	O��o�ͩr�Alȅ��o��)�?�P���/J��(��)>�-��qQ֒7�������q��a$��7�N#&msܪ��/pѱ3���H굪F�H%n�58��G̮��*�'B�87�����%n�p!=ExC���'�'�F�+�,�2���(w�Q���Y�� Y�XO�Y;�2�����dI/#|�%��z�0%%��=J������8��]�@y�? gnd�ns��O���kI�dv�E���E�/%����@���q�L}@N?:D���,lJ�#˩��fh7zC���[��K�1Æ�5��Y��5�UEd��{V �8�f͙��:P�h9_���%\�}����7�E�P�E���E��1D;I�8}��rO�C��\�&�Z������8{3ͭ�M&ވ
 p�����4�BtuP'^
��/�Q���[�$���%��U7��Ĕ����v�����Z���*�\�W�U���gj���=}���D�hR#��E0��fi�ۑ��>5eY���3viܵ�e�����hA�v\z��7���r؇�ҭM�iPP6ֳ}��=����u����!x/�E�`�%��c�<���,G��
7Ŵl3���}S�A�:1��	�p�����_�ð5=߉|Xj�W-G4�Ҧ4�����[�8���UP@����m}M*�Q�CQ�{�nK+hb�M��զ�Z{m���JM�W���1���7����h��PO��)�y�~�6�{�$U��F 3��U_���h �=�������l_G�R*�MF)'<���H�~V��BI��vp�66.�+up�nf�p�y��ˬ�������%��#Ҿ��� *b?0r�p )�ʮ_FCg�^�u�NkRa�lI5�x@�	Ub?)�Y�����𷌌z�|�<04�'�m�r%h?�c�;�_O��Q��I�F��bW��9`&aL�8�S�I)�P��M�~3���Kx����ދ���2���qc��)v���4Z�p�o��I��	�jk���4��V����V6��2@:\WD�5F%�D��o��پM��g�\�!��@�����[�Qxa��F]����/���mA�zl tG[r,?ɳ��h|f�C�f�xgW���tg���	Q�!� ����<�2���
��S�����uʫ�H�1c ��$7ے�]9iJ%��K��x|H��?�u�R��䥏�~�ꄍ������p..�Y�ܬ�ܨpS{�!N����� ^g5K��;U�|0�.~\�p��Y-8/�ة�{^|�1��жٟ�Z:k�2rc���yrS���\�M�A�ǭu��w{ۗ�)���濆���w��Xw�/��}��6�'�Z
��b�!�|��լ8#��;�o7���i��I[�P}����Ę�-���;ɵ��,�E.r���aUț��j���}9$���LZ��N�����Sw�웩N^7+Q�ZrDoo�n&���.G1`��8C�
�v�Rl~Yk���J?:>F JM=߹5���%��'ב�pB�U����V��Q���&3��]M}��L�؁����Ц@q%���v���ߵ�y$Ϥ w� ��?��unin��}�[C�y���a	t³�{�}�^���T�U74L-��9�U#��!`ƕ4:� fPpF����v�N��z$9�;q9���cO����{�m?Z۬.j���Fw�*�6��k ��A�R  ��N�2Ͱmz�����B�?7&&��g�Q7��p�%Q�p��*��۹M�[.ԉ�xKK�s�4����e��".�1* �0A�Yc2�PH(i6D�w�`bQ eZ�:�tb�y9%<�	, �b�����C��+�a���&ղ����;[K�������`����E	�sy֝�w��E��W���������̃VެGG�S��tך��X�����،�����)�U�<��x���~�ݹ�l��{Sj�w�)�ƺ�a���k������y`eQ΁r^��;J��r�2m�慗B�OQ9%$�&Yj���C��̪0�[�E�^l�k��Y���/'�O@mILdw��h�7�܉2���c��_q�������1c����~��#nY�JB��g&jfE�rP+�" bzC�Øp��x]�U��� �I�����gN�@X�5`/9�䊌,�&��>�<p��s�ǆ���zu�k@���9N�v�o��=�	��y�Z�k�.�>Q���+	�R��igF�̚��T�Ǟ	����<D��7w���vUk��ٔ����*�'��'L�.��-�� q[PV���eOǻ�W�q˒0P������sۢ�V�SY�n"�T�N4@�y�M�ܟi��{f�=E�}|��_��#��2����W/4oT���=B�`H�֙�ɚ��JS:Ed�!e�%`��n���q�v\.��p�p��]�l�(��"�J\𘵾V�v�m��g�B5>�w�'�%� ^p
q�nބx��+��>�f������k�Wj��|��j���o��_�ʈ{K`"��vZ�,�[����=*w��Y�R������i���
��[˵��ж����,�"8�s/�(a���M��;�?Zr7(l��U� � 5<��N5�?�Zxn���~Rx�$}I,�OYQ(���8�-�z^��-$�W������0cg���Z�	ȋ�)��R�dA=͸���z������Y�\�+zl���y��8Ϻ�q�=�����6:8m�R��N���`-�J|�����,��!V#>N��Oq�g_�"t�uU���hX7o�m�i�Rr,L��z�->�#8ÀU�#�	6�s���Q69��&��w~�4�~���VC���� "�����y\U��j(�S�����Σ�Z�X�k�O	�!�$�~Q��X5�fѐ���,�4�#u]�1N�.8F=�Пux���|���(��:'�/C��[<�AVĐ!�j����˧��1���:�
�]�}1��L9�?eۼ2K����l�vr:��{��_�3I�p��P���fۼ	O����(a����w��r������̒I|=�����|K���'wJ1OU�#�AT?�^
q.b���\�kr���͸洘�%�Ct3˨��A�|ؕ��`�� �~�Τ$�-�'[
iXS���J;c�wso�H�=�
�w�HKP�~�^:=�!���B��3'�z��G����Oʑ=<!?]`;
�6�������H�&��5U��,/���P�}��մڢ
3V���\[@�e	O��i̝�KBm]�V9�}22�)�u1z��I���B66)X&�ր��1n ���Ph�ĉ��ۘ���BG�AAa��S}}ɯ�*��I��z���C�;i�F�DV�O�	�GV6F�2<��v�����'�/qK�E(�Wኬ��b>��Jbd<���T<�VJJJis]]p�R���SM����3�rW�����BF���7��!�����x����!w@=l̺�㮌c��*3��ڂ�L�/��"U`�*_�!��?��^�S?�z���I�^E��[�ןb��R�G#��ݎ�]���z@�������]ϣ[Cگ,��j=���j����4ݗ=��ڱ��Tu�:$sy�ab���0d��1�L ����G����5�>9�iزiK�VFQ�f���u��?FSS���X^s��Ja:���?QY�����]ǁ�%��[����n�t���>cd�n���5��e�#n�{~co׼�X�LJ���%��2���W�`�ee*���K0Ȭ��RX}	y�q��/����(���L.,~�{�r�*�Ţh�H@n=w�-�˄M�8�sũ
�Z�1����sqw��5?�mVYuz>��7P\�?5�*l���R���"�<=�j�"���3��ՙ����-$ ����I�7n���b���1g$���i�����9���L/��q�#������&�FFJz3�U(SR�S��y�.��@*�'Q1���X]�./��f*�����'��$::��Q}kY�u!>K��~�K��z6x��0晀k�˻:ݴ�+#x+A�`w7�s�dm��q/ɵ����\�ig �ִZ�$���H)���Hd�g��u��#�.����[S"��u:�
8��k5Б�~�(4�}��iM#�����32y5r�`K���\c���׍���g,�d���qJ(�HDKR�Wuk�WY�
�ym�fg�ؒǽ2SI)W����qȮԒ����+�ϡ�36ZB�!B��V�	�(�dϓ�S�,�g�����g�Ih�Hx��Ȟ��|�b��.8x������+\b��O�	������_�K9f�Ð��n��T-�w�s�Ǻ�奯O�F�e3^�����"X���/)7�z
l�50v^���f� �T��剡��O�Z�'�jJڊM�6Q�PK   6f�X�Ƚ׌  �  /   images/9185dcb2-65ea-4de0-8d42-42cedb1b5634.png�x��PNG

   IHDR   d   -   X���   	pHYs  �  ��iTS   tEXtSoftware www.inkscape.org��<  IDATx��\�o��ݙ�����uڗ��!Q�Bp�D"��h(U�$B�F_���?�C�JM�!-�А�J�(�U(I��E�|�^$k�w��u{�ݝ���?���gM|}?~3���眹3'֎_�A`$�M!p�8	Q����~��Ql18���gv`��ű�K�Vr���x�p�z�3���rW�y�4�0Ɲ��t��=�r�Ҙ�xq�!4q]&��:׸:/s����Թn�?V̕%�p���:�+3xg�X�@?��Ⱥ�qO�W�t�G�����X�ѳo���Ij��;m�I�Ae�ŰĠaä���	.���'�eV�	C	��h�*��2�z�=.�q�k��I�%WZ�A�KD����rB����'H)��8�{?J����>�9���v�4�'���~��.��7�'`��9F+ o	�'�!p��/e��!i{?�CP����Ij�Ҹ<즺aj;C}��Ǘsݥ��N\₱�ߧ�$ސK�\��G��	y��s���׸��s��%\�I��,� ^�cg���CT���;s���/��e����2f�f�}x;����Q���r�����2	��b�\͘�#���-��pb�w��u6�S��;92���&�}�5L|�,�a��ʚ�K��D1p�eM�H��ugDq�ߣ�[5.W�z�D
!����	q��MB\s%��Zs9ߦ{�/�$��b	ӓ9����M%wk|ao��3�=�)㭱�I��4Me����K�_�%?�q�<��5'��-����Ү_���W��:�of?�˸S@�w�ۻ��~Ϋ�1\��K�
�^=e4��"������W]�r�\�ո�k��書��հÛ�����$����ǰS6�}�������>��ذ�)���Ty�"��])����ZMtXT^��s�V>�q�<C%C�u�2�~󘫕���M5�;s���R^����D����}�s_!�.I��VH����k!�){a���2��0ڔ[���̵��`@��XxL�zp�f�S�7B��"s���q�<σ���ҿ�P��J��h��Ȝ���g.����U�^}Qx��t:��C�Z%�d)�jдЛ�s�1�J!�H F����R�����Ӓ뺈q��U!�M�#���c��"(�Bt��]R*��V }�����H'��t��Q!���xUH~&a�����!١;غ5 CG�4�O4䏱z��אi4)D�Ζ)�L�8:$�U�vQ������:�Gx��x�.��~���n#���q�EA/W�W�H��s��������/�]]T<���}t��.��j�G�E��WX�_�|BE�
���Y�0��/-S���F�]̓����@�1����n���~k��j�ل�C�ޠهđ��CW�c�+��+���\�B��T����8���u<6:.��aYC[q��Z]C�r��X	�z�Z�Z!�Fcr=�/��Ut���q�@�\Ѱ���\�d�\���r�r>jp������!�=w��B��B����`t{c��	��겻�GA��lZ��v}�m��_�Z��v�qb����/�^�B(JKO���'a��iw4���������~zHي+ڮ���E�S>��W󉞻�S*;e�d��vr�-�+�hVXG���f䫊u�S�#�J��Uj�pc��mw|}���l� i�!�x_~=����oܺ*�5��S������q�8N��\����MW;t}c844��'G5���!����}yB����a9F{(?"�_�$9�c�3TC!���
)|�B�O����ؗ��0�W&�RxT�R����s%v�iѥ)��	^�U��=+���0-zJ(���/����R	o|�6��}� �3n�����=zw�G�X�ξ���z0;���<w����4^y� Ο��R�¬����i�C�8��y,U�0��UI�c��W�1��u�Q��\�����p�{`�OO�0Br��V�u�0���\�=�r�9=�Va2^��ͅ	!�sZ4+���w�n������ة�jep��!b�~?�7�՟�{PiѤ ��?�(�*��    IEND�B`�PK   vb�XT�7Pb #y /   images/c2d54090-2fd1-4cc2-9c7d-28b872c3ce05.png�{e@T]�6J)ݨH�C�J( �0�t�tKJH(�)�=t�ҝC+��Pߙ�~������~�g��g�u]+�Zs���(�'�{����A(+#���q��0��a�����o1J�n�,$%00ʣ�?b�:��8b`�9���[0�w���˖��Pw3؁c�QL���a��♜3��b���<���U�n}��G~XX^��ßP��5H��m����H��I�O����O]�����[4Å�]/�V�E/���[�3�Z�ۋ X�"�����ạ�l_�q���sC��פֿ��y�X�K3�UF�gYs=���}���;fS���Ǡ��.��Rŷܕ���r�s~᩸*��q��]������2��ivh�����Δ5�hg��#�SUut�L�?
�mC\9�!Cϸ�A����#�;�
gx$��Q�WnW}�A����%m���e�������_<v(���B�D�9�t+�̋��B�'�+��
�X��*�{^��V��IΣ���R.ޟEnzޡ��$�<{?�p��'�����cWl F���x�Ep�\�)�y"N����gy�����A���hv/jK~g��"�	��K������������-���������nX���j����؎5���BQ���;Y��i��wvL�̂�R=�:Q������
~?^�$Ɠ7�r4nSjEk)�7��7'�L��<E��ţ�)/|!�ٙ-,��y��J����S\S3���wh���(ݓiM+�VmU��V@�D��фZg|�Je�,��+FY]�%�!װ?�;l*w�\�k�G�h��2E�!�B�6�����3�v�z����`�sϱ��	���D�ް}{]Jx�;��SS���p��Wݖa+���o!r��3�-u��C ����y�Z�96qžW>,��H��5���㻫�A�?=?�)�����J���Mգ���}����c㰋��B�i=o����N��Mrg��M�O�W�F�t����}F�|���l&D37�Ns$�[����R`��Q��a
��4���p�ӥ�Jxxû2�[��u������F�X
����M��7G�s�#���r}�9$!�=hg������6��\�+v礕΅��ml�[}a�"i���Yy�$����هr7 ��.ڼ�<˯�C}�u]U�fK`�Bp��Xi�8�Ĥom"x����f��o�_ʪ�%���kR�s�.Û�7�`��?�+󕭛OvX̬	���C���\8�Ҽ�A��V:�ӭ�(�
��-���� ᾵1�E5Cc�ȿ�od��pJ�)�\{:!�/����s�Zn�;��Ҥ"�h&�I;nܹ���~o�o�qi���$y�ؾ����%�#v����h6S,��	��&<���	�1���L�ޏQ��#��6��O5��&y�w�vI�r&��M���O�J'�BPf�/8_ld?W��	1�il���2��\E���^ʰ�r�bD"�R�A*�ߡC�d���$����վ����R^;!,��ZmdO"�XE
10W���F�s[�\��Tĵ��_��~>?`�]_����ǀ4熿o�]�j�eV��RC�4K��}aʈ�K;&6�@�@�ܽ
a��1��9x��RW����t�����Q0 [��8���˃��8�b�Q�Rs��VG�眆��Jmk��rw�-��I�U�U��-�]{�Z��ߖ߽>ť�,�(��Zt����ȏ7�t�Ɯ��B�|	�1j�=����],�{�"v��֊iLH�f},��c?��`�Ą���|�h����]R�$}de4em����ZqqR�)���A%x�Az��‏g���|H�����	����NY]n[�N'�5Ce������HoN*=a��1ʛ���X�$P���\깍b�&I=)_YM��0��]YT[׺�_5�a�����i>;��>U�6ts�P�~s��[�<ͨ�꨾<GC�3��� �X���r��<>H_�}q�͡��?"*�7bJ��ߔQxŋetыy���n�SK��З��J5[^{ͅL��"��I��
}D��|��K> ��2p�d;~$i�v*~vs�X�NA��͠qǋ�I΀�2�/h�1E�(i��������yL���m$�w1Xt�u�2"��f�f��J[FQ�}��as��S��n�S����h�9�W�%���ʢJɄXx*�S�G7/�.x��٧+�|Ҥ\�l��ֈ���W(��%n����5���{�o<7�؅d�2��0��W���(G���jH 2ਓce�BG!���'&��^��{���O���Tw�*_�m*�@QK���\gl�q_�̮2M�t��=�JRe��9Y�I�ʨ| ����%�l��ٜ:�B�v���c<2��O�I,DD�hGC|�N
M��׳��G�`�t*^;��K��9E�%��\��(��qЧ��ޑt�	����1-nG;0dwMq��Հ��A��������8����,G����yi>P.7�O-��q]Y%K��� �&D�nm�]ĳ���}�S�o2����.���� ��� ���"�������'��y�BoN�r��0�~ٯ���,�����z��Z��ԧ��d�T�c�8۳���>�e�����w�(��:�1��0��"p�)��d��4�צ�$5�W�K 8I<ea����Lǳ6j��'#ѿ{3���A̋ [a�r�*��<d�=r�-�&5>��x�ܢ��!�!:[���H������G�l�V}�=Jo�0�]t҄?#��x~�7
����|r���z{�����1��Z����ܹZ}���6~\@�dXsg�~�W�>l[H�d�GP�	���͞�s���e��2gL;<2j��R(í��ӄ�K��o>�p�0c�Om,�7�E��h��6��1��|��O�;h���[ntt�wU��(sp���*0�~�2����ܭ*{�N���Υ(�qj��8^7�zr��<O��߲|����#��Y�2�$Ov�R�w�i��-���keozu2ht�a�`ML���;��_���r�vG+�'��XE�pM��x�E MB�yv�t�j��Z�#�L=���jj%ZlG�!lw�'d����S	%*}ƞ�(��D�
�[7����X�9��:NJ?M&���I�}r��� ��8��5-D[�"N�Q�jIrz"�K-9x����/5�>1���,{�5}��Ԕ�,��|��|1��Ρ�:˥���#�U�H3���:�%r�n�1�"`t���}�]��ˌl�$쳚���4���.]���d$���	_�Äw�����!�X�7���P ��xX�Tef��c=�"�o0����}d
	5Ƞ!}'f�Ut)����@��'�xd��|K� (��� n�.��j��0�����w�JkƦfO����/����R�S���������/�4�؍��⑰��[�y�������Ə8�ﱊy(\��_�$���q|1���N�� �G/�4l�o��u�R�T��P�j~�IhYzq(;��$2%זs�G��N���E�T���QG}UM����z7�m�G���8h���t(�sB#�;�{��l�m��eNS,��Q��?4s"y/Z��7�s9�)�%�t�M��N���k� ��5c7�\k.�8�2�Ac�~]�K]������l�����[�b���!k���g.��e���ZY��$���E�'آ0�[3E�m� �9Yd C�u��K�uhwɂ�z�r�t{?�+��h�z���:�|��1N?���}r�X�F0!f���kU���AD����x�y��}@u7���3$�w�KZO�R��|6��� A�?/,�d �20R���l���� ��O���5$Z�Ͻ��6��4D7��8�6@��e����Ӻ���m��I����GIl��$f%9tY��*/^��]�j0�ׁヒ�ѥ�GM�=�k�I���>ɗ_�v&��X�R	 u[ӝgc� Y���g!J�v���b2 ����[�7��oYpp'$&/��^.�T��\��막�}o,��)P����1>���9U�0j�Z��ZF����
��85_���֬�^!.~�w�+�E�PnZM|㼷�۽�OhS�}��ߕ9Ӽ:���[�o{Y�W��Q���N�W����/t��,X�T�Aݖ��@��[�UuD���u�7*F�.���IQ�n��q�Q�Ua�4�$vZs)@���*�hm��B��݅~����-�KZ��ƨ�vR�UG�	��>C�V;]��ԙj��rӆ�H���Ȁ��*n��(�T0���9�,F�)��I���9����7t<y���f�]�,(SJ��2�F<�ss��d�|�Klv�s�t���|�xB���M�g�'&��G��sf���j�k,���{���WȆ6���H��乕?����G��1�$�6��s'�����o���m��ZB�3��*�aUU��NՈ��/�֗�9�qyW�ɢ���d*�M)��WO���wc�]4�}'����w'�Lܞ�-�]�٧4��_ c`��&j�a�q��9W�.�E��7puB���	�(�FD��+�E��_�L(���QT�;��Z�Y+ѕ����vF��z\>����mwZ$�\�l�7�ۣ��-�Wڅ�?&������^ �{2���7;ۥ߫,��L_7��/)gٴ'�b�H�����N��zµ�"gm�01�yE���C�q��Q�?��<uO���'i]���J��sk[��AD��W�Nh*xi7����|řn���lua����aV��b���
���J�2�����A|�`3��s����*�{�
�m\�tX4�,!����<�?����~���a���^�]]r�ɆR�}�&�%\�c3
�`�7>��ܙ�����+z��ڼ�/)h'T�~��7&'�M-u���b�8���L0@��#�m�� .�� �&���<d+�2|3�xaj��ә;�`�y�>w"N���U�f�^�w�D���D.������|v�� VZ�����4�@o\�8�-u-|}�#���I�ދF�	[u���P����ū�A���B��)�S�@$ѝM�ً-H����A�uZ�
��LU�T?R��"�)�gZ��n�.R=_^lJ���℅�MQ�6ޚ�+���R���:�@� ��ɩk�4�R/|�X+�2���Ziط<�a��F[.S�VW��+;�������2�	�����ʽc)J��o�k1�(��)݄;h�*�h�w�f���oF݄��.bj�˒��̿�$��/�99u/��[&s���Uvښ�Gʶ��Q>B$ �уuW��-ӿU�0"�el\��*��l� ��]S����Oa�%L�JRU��o|V�wl�"5��$́/Dk:��W�Հ*@����?���r�V��'6'iZ��� _㣠�|��mſ��oX��2����<�n\M�A���OE���G"�4��H@���yn�n��]�ڌ����M�� �@��1�^ks��@�$w��!#��y^�)�{L�)�=��J&��O��qVl|Y�HS#�x娽aT]�^�y�Y�ii�zv1�P}v^+��
7��/ԛܟ��	T�y2�SA1v�"	m6�J���h��E��ώRs��$Q�Bl���;/�yn��������1ub;���i�]�����h)��D������]�rg0��u�e�m�9�~w{�����M�#� 0@�K��Jl|���<�Ӛ0	Ӄ!]��6�v�Iyl�$��1D�6��S)/97��F&?B��B.�U֡�)�<��>�F�j'L�Kk������p�:���v��b\u����֐GV)n��`[�e��o�U2A{w⸽�b�n\��,&.o�DHf9�P���u���/̻���^����s�^����mO��NF�}�K�\���l��j���kB|!��Y��:�It���B]��_�k�L���#Q�(���]�3/5��
���0&6�P��]	?	���;��v�0{z���la՟�K��z����C��lLk�PMg��I�؉�ʡ��HEˌ.��/2%�F�b����b��Ǉ���+G�2$�Z�_R�.Y��S�U^�^��  ����Ԫn�6�\�`��K-���G���r79���)<�E���n�Q94Y�0�������i~��$M�Y�E���J4�b3ZM����Q�����pѫ5w�)r�t���.Kg�M%�[]��\�.�y���֔ւ��w�ᕣ�<�4�ݗI���R�v;0q�k�ڒ}R=�V#TM��W'}<b64�F�=�����n�a�����;�N���2䱿U�X�����Jv�I\�5���tE'(�V�R���y{�J��ދ	�7�v�����X��d&<B�5�҉�e���%��X8�6]�t�Й�A�_eQ�c)d�.�$L�
�n�x���k6���:�wN���(�-��vt�R�+�� ��:�#�&�-������+����=����O�:�ж���.��}��x�s�HR���qiKN��^�Y�q&H�ݝ���f��U�д������T��ѓ�	l�7	�Co�Q��
�o�|�$�K��}�),
�����������Ì�]m0�ɠ,m�g��Mғ���]���qy����S�d����ކ��D^;(�!e��͇��RO�vf9>~qp��C��3eu���Bٖ��FX�H����d����3�6俓�Ҙ�11n}�ɳ�sA���m)�_���{��j�W��=V�@�ji|S}�9�SK�&��N��vx�Fw�c�p7�EC�CLG�"~mw�>��0�O�������WB��z�_��Tۂ��N�Nͻ0ǜ⛎p���5����������)j9�7��]_�{^_���掝�4F���?.�}	�3�F`%?��~�F��������*��(�����������~���N����&�~+R� k'�>�nǛ=�:�pY�X-m��ڋ���=T���Y8���)��B��
�������Wt��k#�J���4{�p��=5��{&�)ee;�v5\USjh���h�.�5�n8:�w�WV�PL>����@�߫�����h�]�����s�0�.�ٛ�-�@�I��7��޵%��9�;�ӜY٭P�Ҏ��ˣ��ѓ�t����ҁ��\ц��s��]+c%�G�F�K��Db�1=Sb��rt���@�,ez�7l8ߢ��%��h���鼛��ĉ�@ކ���#B|k8�t��!	�.=��A��"�w�"�#ϐ��_R���j�a�^poX���}|�E�)iD�n�b�u6PO_�M�
1mXl9c��MX�%�B�P�)O���!^[q(į[�<`NLOW��?�
X������2Bo��&�8
�ϙs�kAR�����_[�Y�^+�;�[��	���e{��sg;�7w23s�	���R�P:Zu�X�m�rgϬ�[����
z2�
,M*�`XV
D�p���u�Y%�5,��ct�?��.��?yK��1#�D2��}�N,]�����m-��ʂ� �������סBf6Nx��%,�P-�˴i���̽�b�%��� 1qg�i7�SႸW���q��H\_Y���������!�ޥ)zY]f>�@���c+�C�ݖ��9+��B�N��(��Y]Ț��J����=D4�y��pR2�aly*o1v4�"�d��������dIuc'��P���b'% þ:`�ƍ!*X���<z�pyoxa�YۏO���[L��<&��u�"�� ���[��{��
�<+���kq���Ғ�+V�<���,��j�������ٻ�MYSu�ݬ���Tvښ�(h��ʇ�	Ѕ�3 0�j9g��Vo���X�5Ȳ�XB$�63�8g�ZJNc ɔB\v���t�k�7�� 
"�8F��wk}R˫P���;/4"�}n�Rj��88+�!$,oJ�s��"�ׇ��V����� �@u��9���m���<l(��¬�H�ޑ=���I������������JY+�&`t�}R-�����0
6���}�fV݄��F4K�%�^��$��YoL2y��k��Yh�����V3�RE�Dd�Ul��d QH���E,��|�R��:�d��/���d>^����$A��Z!=l;b���]�r^�z����Z�lv~����D�h�c�xK�+`cF&S��J�0�f�|�}�a��F�;������@ ��N�=���I#X�'���̒�|D��(���E�i|�J�́b�H�|Կ�;_�� �%�|m=�k�����Q
���1��$=�/e�3�p�d @ 1_���V\��D������P�0�Y�<X�6�9|����dS�����2u��>y�X���t�`j�{�
,*�G�V
�	_3�\���ְv��($�߻��4�2H����	�����4��4��`ù��	R���`�~\���XT_���O~63R/��'w]��˚���Fh�����jI�@�3����n�e�.�=����-�U��n|�"�%QO��$�gt�<Ȍa�%ڭ��|��[�Z�1��>+��\K�q!I��.�֟����K���3Rʱ+�|��o[;�/�o�aΡI�K��4��\�G��?�Y�"�Se��sm���-ѻ�϶��u���(KEa;���`T��a����z�6S ��˞и�0b�l5�]w�����h?���?��\=⪕��Q�Y2���Y��TYgⶴQ�һ'F�w�K2�ˆ�� �]��l���g��EI��G��2[�����P����'x����[X1� ��E�K�O��ā/֫n[4�u��{�	�Ho ^$�L��p����Uq�V�e��!����Oie��.(���d��2�꭛�H�-�5����Y��!W�
B˖�#�8��&��ބi$[a�8�˪����[��܆���~q��F�޽���N�7I�0?˲Y���u����̂�_�p��g�J��@�����Gܥ�"o�X}v�<!����c9s�Y�8��v��6�ib!�_���Q�`�gH�h�_)5�Gg��O�xkn?*H-[Щ��fe�̻��z��k93[���Vc9���V�Fc�����@Hp0z�(<����q����q�����-��Q�X}��>�(��s��hY��IHuxq���uͅL�"	�u�ײ�*�� �o]e�����6��]��1�b������]�X�=vPg���H�Ɔݐ�O���#[�ޝu����e^�C	��������:�3��未�A4����,�M�-)�[Q�K�����Z�����֕��Vkc`6����txǎU�QT#�@�l��A I�Wc�Q��1�́'��5�zn�_�Ћ��i^���|�6GE� ����iC�-���Kܐ�zJ=H���+������5�������� �h��K�Y~�����Z��T���}x�H,	����q���2N~`T�+mc����í���3�J$��[�J��w3Cpa��E^��/� >1O	��iuN�>��h𲕄��Σ���wh�u�k:��?����r�����SxP{���wry꫷����s{/��*�#*�°l�W�jYf��y� ��&u��>H}��$�'�����L�#��9�'�d'9t�Ckm���ڶ��I� �A%D�<��_�i��)B��c@�(W�^�&D�[�+h��K���L�<r��Ӯ�����a��A/@|n�f�F�IK�o{K����zőqnt�]��G����x��|����w�Ó��yur������9'`�;����!��:����y<�M
���e��:Yh�؍���� ����)����%�O�&�Z�dc��y��sw<�A��w��>mؗm0z�)#2�Op���Sb��<-t�3�(��Fv�g�����.��O����`�
O<j��_K�����!��0�1L?��G�c�t���m�~iD?cw�o�g����Ȗ�M'�Q� `.#�=���K8�DMr��>4��$$��Wa]v�oܟ�0*7��j��^.+�s��[k�p͗��m^�l8�}0�]���Ċ�|ù�[�5���(�{�e��@��W�n0vʈ�t���5�I�� �^�eY���8�t�_A_K�q���Ns�\�L�J�Ƣ V� ����3O��2۳�{#�IU2̒�cp���}7�vrx�uW��ٳo�Ŭ��y��cD�ᝥ/Ӂ�ť@c{����#��	�%��#e�~�NBm��@��z����t�\
@���Lҷ���ϻ����Z�я�x);>;�m�~���"����g؛����a����F�����rL� �jl�.xU��u����v�T'����o!}%�҄C�.x���E��u��z���DB�tPץ�s:�*0�_��^x�)��3��������@�^�\�X�eH��UD]��$��Z��T�8)����F75yR)]�Ac���ڜ~�j�]Ci.@�ȟ =Շ�jjzwBY�G=ig����8�@���s���A�/�gJL�1��h���n-�7*���t��		�с<�|�5?��	�PF/���������J�=�+�g;=�Y��3tД��ؼ��Ǯ�9�QQ��� S��/�E����N)������(�����N���T��2�i���g%��ƙ2�).��e�Co@\o(�ZJo�D��h�"��9&`�"��-�ƙ{2$&V�=�Y�Nn�K��Š&�A���S`��I�W���6����YV�E�E���Í�ʍ���_�����������P��ů�&C�-��'�F�`��턆�)UG`gh�苍<&���V�/�n��V��&!}�[|���kNӺ|�y�����ӄ���k�y���m�_�Z#FqLȃ+a�|N W��	 B����������p�����.���|��B��sNF:P�z�Nɢv����ftf�Z�7eL?NDwp�sN�Ձ9\^b��`�\pR��ܐry��%�mLRh�^N��يc;��W�F�!��1ږ��;k~�{���}w�WuT]�E(��4m�Ru�F�E����՜Tq��v�v����Z��K�CJ���0� ���r�j&,pD,�W�n��&��<t?�����2q_��eF�b߽�b�+B)����?Oc��E+��r�����0�x~�XP��/U)�ra�X"����De �Y����Iy��j&PL��N~~�`�/3�R��.~o6����Z�gc�D�WQ��V#p�_�8�ZC��UBS���M�
Z=r�`�b	�m�
��{���}P���$ �w���� )Uֶ�H}]��!�H�y��IF�c�{�H<�'��VvQ~��� ��`ӍڹV�Zn3-\�Y�� ��<�C�w9�ps���Q���AP��
��d��������>Ns���Em�&�}RJ�hn����B���@�lw���8^"��"
���B`%�U�;�H�16g�u�q��`�TA��%�<��P5)Ąb�����3��U>~E\�˂&�T�L���x��%z3���m��$P�UZ���^�+�J޲t)D� m����,g&����>��E "f��IE"���j:�=�a����s��Q������!v���.s3���Al���)iQ����1a��r*2��g���'::�����93[K6��99ubo�~��Sh��O�k&�0b��|��0j����y[M�E-H ����s��fhp2���)r�9�z��4)��n���4j���-)���n=��ߙ`&���Ee�]��b�Ў�HS�4��_����g@ƅ��Ĉ��i��=/xP;*U
�w@�Ȏ,=�!�%��u��u��l�����ļ�]��o��3f�HEe�E��_�Fmݙ�<�Χ�hv�G�-h�d�;l�mL��O3���
1ѱ���"iFs���O�}�O���<��55��kj�r�Zb~�ff�VN0?��� ��% ,	�l=��VZ!~�ς/���k�z��V+>�Q���$����m��-�le�<$:�0U ~t\���3�4'�>�����y�TQ��'��>a5�j��x�����*63%�?���)��;,�"d�j�s�!���2���qtrK���%��M�K��jr�8槓=��)�P���.�I%��O�1�J�"��EOt��s (�5���v�EǢӮM��e��Ȟ���#$$�(ڿ��*����eX8`tg+Iɟ�Tr\xBe�F1z� XX���^:�l4����pOK�~���x���c^��А��ܕ��?{����TA���>���q���	G��l{�@W�L����V:�,As�jkÃQY�r�?��Z��G=�����
�V˭�4RM�jU��v;�:8:���wk�)G=�c�L�ɘ!/�E�ڋ%u�F.�oĢ��@A�r�S�n�T�CS�UiD]�b=ϣ׏�R�i��� �7ռ��:e�*'�J&P�yhI� �"T�ߊ�c�}��Mb2%PJ�?.f���Ph��u_�g�K	�)DD"L�O^.��e���;G:�SH"�koŴ��DaTHI]=ҧ��#��:��O����%�~�+dAV��-A!�|�"˿Y�O?5�!�K�D����2�ۡ6(�K�]�����	4��;�G}�43�\�Fȯ���E�2�����f���E$�е�����'w���Pn�ߪv�B�y
הc�pmI`���H�h!�R�Qr}�������B��Z6�Bʙo����f��	��H��D�5j�b?��>�5ÁON��q���������}\�c�����Q�>}о��4r/u�ֆ>I�CT��*��6�uϐ�F,*l!#����@+�Ļ5f>���U�yY�~�v�J,[w��w/$�n�ɫ�	T��[_�I�d�7lFl��̩�.�#O�jR:�$���S;]~A�s6��r ��ý<PG+<;�szdr�;��A�s�4�/$ԏ׿�/�7'��l׌�>^�V4@8+s�L!�� ��+��ce�S��h
au�4�a����Z3���v��E�Fͭ������?���/�OIN���I����[В}�<NjM�-)���Yw#E�KW�Ѓ����K�Vo/I����葈��RJX�?Gn�z��AIo��� �������aG�-�i˥	��`'D�m��[v���E�c��;z:~6�dǦ�"Ɂ����[m�b�U��C�������80r��������b�M}�9�����|ϝ��evn�>�bJ��R^�#
�P$�Qװ�Zc�,����͐;����t�Cmi;HB�>�͛%���psD2��8�����{J��� ��c��R,M�����Y
%r|���B���k�$c�u����diz��X`޽�)�VA�GI�� r�!ݰ	
[:�|q��7}'$�H7�t}z�x�˟r�p��(��d/��wWP-�i{R}�F{jd�{T��f�d[��_o��bMk�JkR}�4-�Xo!c�β�/� ��e<����J}.2A�V�+��!/0�9a��Ht�1$��m(��u@y	G��<4\6����׏���)v5����:^-�K}J�(��"�i.\��*f�/P����_���wO�&�	[$��/�a��L;� N܄':g�O�ca6ؽRK�T��7̪Ѽ�I�,�w��L܀f�>����nǕ���%��+�1�@�r;:|�@�P����z��F΋״�:#5��MJ���:���ǵ������I�Qt.��U�������Û�I�˯b��mH>�>$�:�2:p{������RUe�װ5��� B�L�g����̹���d��q~�b����&Q����Xĵ4[�5��#�#�d5y�cEƩ	�P�G�{`�8�aO��X���t7���kμ�Y�t	6h�o4�lCG�����#����{ �Ɣ:�m2~��+�Z�y4��t>�꫞b<f��ϕ�9x�h��\�c�A��0�o���Jc�(�џ_�]�o�{&���y�<�����v�݅Y�P	l%t�U�!�K;���($�hS4�͸z����~K �J�;�N��#Lo�����S�����Z��b\|�ф�%g�B��%͕Ҍ/�&���=�E�_-�]j>$�x��zx���B��޻�������5��WM�	4p���/,��S�l,��E���@��^?`��=3��L|fC��u�C/ɞŬ��q<E�{�|�y6I�"Q�{	�-wXs�z'�5�<؎���[j�vq����bu��kS��I�X09^������Ϡ1�)�Q���q�����}���X�p�O3E���0~]�C��~��;�	���zb��3�9re�YI��{�˺��Չ�n�U�Т��
OX�Bf�V����+j��#�Ҙ�{F��I���&�h<�=.���p�8�bat&7Ԗ�I|�f)����a�d�p���7�螖�YW�sN\qHN�@,з}%���<v^��t.�^�ZuF����&�9,�q%n�R�a0�Y-�%�Z�����=	 E� 7��W�*A�7K�.D[<\�XT�J퇉���z$����d�U��3�G���ת��P1f6eAH��tPO���t?i��H�'y��L|��ƀ*�nԵM��4,�܁�v�$zӿ����j�r|ojS^��?T'b��D�c�o�w��vL(�9@�&��\W��JA�H7�V����bje�FN��/��!��+fN�$O,e=2\�K逯�򦆵o},�r��Nbt�I���Kk�n
4Eq�#�b��N�#���=��mK�P<�I�I�<JX̠�t� C�i�J���[�.m��(��|(9�68�t��{-<x�*���S�������-�2#.�2�;�R���/!��YC3��'�`��_�����+�1�V���f��w���!�/}�EeWG��������:Z��=��}���dbl(�N��y)V��5yk\��3�yO�6K��-d��N����-���F�d��\��Z�����5�����ɝlx?ewn��CAk����h��������4�g~��s�^G�N<�&��A<���d��F����h��Զ��~���"k9֑��Jo���+TF�U9~�J�O�6]с���l�A�ڼ�$�f���
ȤW��_��\BخF��}A���G�3��ZBlF�*&��� i�=�'�{�h���Y� e��X�s��a�;[V���_�K���H�wn�y2Q��I��x,*��(�f�mM��O��U��h���Ч��$�@���Þ(���x���7��^9��}��}���o@6��Oe�\)�J��z��v:��OK���Ť�X�"L�'��`��5#�瓺�cq��w~r�C�V̑ď��"l���ԁ���x�O�#�zUv��_I�.� �$��c��������0�0R�ǎ�!�J��3��`�`�nD�O���^F����%44��M�"d]�a��rLiv�Et��.TX���O��碤E��]�w�t��kd[8$�)�	l5���O�`���
����1���GY��G�|P󟗃�de�#(���v呼~�e�hݸ8���1��C��:~���۪��~�s�րU�'a�@�V�l���s	A�\�����`P>��^j�m�]�l�����勖��ٹ	��>(ΈR���R�����#w�Ub`4~g��UC��l@��VW�!�<�HPf��<jsa����7�5�t�T+����2n���rÍ�A�ї>�鞯5�Z�����z����k�=�5Vy�@�T�B��#�������p��';`����$���y���j���UH���P|?\��al��ъ�c<������z0�khN�k�,6�KL�`+�=No��l�C��8�8 ��"�OLhu�k^{'|d�2��6'f���hbq�	<:�����D�"�D[Շ�6�ַ;J2�Z	��?�=�g+`�_pu.�+(�U��9�ǔ��N|ݺJ�0?�7|sM�?���_�h��tI���U�ܥp
u��LY���3�9ˢؠw�YK�COf�p�%b������H*�4�bo�wlf��� ����~&{�9�������֋Æ�4�Т�|����'�{��:�k|��:�F�R~�c��냩K/T�2~S[�
>�;$'bhӅ:o�͊q����n�l�C�����â��w��
����]�1��i9l��*#�G\��W1̙k�닾j�q���6=_l����'(��d@����ކr
���?�������V���1�/�9X��G-'�8�q*��I�©�b��������b	�����]I5;�#���Zӆ�fP&�Ւ�!1�������Y)�>���\$Ӑ{,��;��[����p�]h����i^����3�0��c
'����;��v�<��]�`�������/<�Ҙƿ��_����~'�v9Pk�+:Vԁ�	�zI���R�qT�L�bF�UQOt=�Q��i%�g�
ǟD9�l?Uk��U]4�?��u�Y�ZhL�&#3{�mβ�x���??'���Р���8d9A41(�)��l�^ŧM�T�Z�x}�_�����tH��@1�'��"�����,�D#'�~�8� �yj�'��A��e��7wVgj|0�Br~��x(�P���y�?��:(�g[�!w<X�����w'�����]	���]<08��~����[�����j������z����{z��;OV�����(�K�?��L �Jpҽ�S�xs\�T�"1��>�FM�ɩߑ{���#���S^o�x~J�e,�yy�i^\l����CF��
���&
P�a�$Ю��]>�D�	[���ֺL'>�Q����s�uؔ�9H��~l���k�n��T����oC����>K��:O��#��\Q�%.ȴ���1 Q4,�%I�����P赦��[�c�n��,Hl��-��]˗���䙋�9� P��2p��10��t��w�TF;�*?�����_��g�A'0�i��~�g(0�:��Z
*
�aQ�{����,=�Z��/Vɍ��mé��J��=D�㐱����hK�L��Y����1�
7���T�,�B�� ��u^U�����0��N��!x)��Є�!Y�A(&�'�	����咹/�|w�˗�~��Ľ��f�g$��X`T4=��y�B�"���Gr~t-f$֤�W	�j���}i�&!�@w�sP�6�^&D��&1�ֻ��S�Z��Ej�n�`�-"ғW@��,�a����{]*���'���%��k*��l$��d�,�lFn�Y��������Ś2�D��4���
����7�w76�A0��e���2S��"Et�a5���  ��ʪ޳�հH��?Z��c}^�}��A]4��WXG_;��[x���oB6�H�f�z��A�]�9�.�p���-�lJ;}C��2ʌ(��As�_�� >�a-;��{ׯz����R�5�{Ld]~I��Vw��������c�hJ+'�w�g�DLn�����l�\A	sv,�6~aV�!�����S�{c��:�n\�_<�����+"eE�V�%����ϮQY~@L��:���Հbj���U
-m�f��.�Tk�p���왔ȘX��.ڻ�
Yɕ�Dל��腹i�V��qF>�p+��T�D'[houy��N�gʠ���zH旡S���f�	�N�yw2�(��H E�Ԟ�@�uYk�$kZ@[%�c�ț��DX
�~���Cd��~�L~{W*?�tlx��L�j���uW�����,h2�2��?nz<KF���.d*{��#xHmюWjWsC*�A�hwQ���L�,�n�r*���{ݦT�Y*-^��f��K[Je��	L�ϲ7����K��=K�t�d4�Z��1�B�⊱-�]�1����Kt��C����(�]f�]��f?���xe�5kIa�C��C��s���������
S�LS2l��U��T��,%���-z��-��"�o��;W�k�Z��i\�5lb�(��J,
�ĄZ1�.>R������7^ݗ���Q4�����66U`�d�Z�K��f�kD���� �ɐ�?�`iʜ\l����@�'�}�0^^�/?CZ���a�=�uy�;w�C$�7�G��e��4�T/F/�F����A�mxq�%{2O�D�(�OA®����m��ɠp���N�la�}���P�=�n���(zF��;؞Ŵ�bxuG����52��	�EC��_��C,����C���vP]�v]Z3�gKT7����l�X�*����.r�����"�͝]�m�e���^���C����5G>�-�H�eܷ"i%M�0�x['�hL� p�VY1���2��e��:=��� �S�4��{�o�0����1����B�=L�ː��c�X �*�%�4�%P<�������Q�,�o1��¹$i�&����Eܡ�!Ic�j_0��?��r�z��{�YJ#$N��p�~|@�+�
�Ra�iG������y������tx�c"��� �c�s�u���xfչa��n&��;D�*5���q��	���M�",���g�?�z�,i.�uW�Y��#s���P�p�Q�V�U�C.�q�o��;N�����O"���M�26�Cw�sn�]k�X�
��-I͉�D���·%@�5C���)���"P�µ8��=�>�˫4L�4�CC%y�83}�|>�S��Cڦ��<��L��	8�jw�N�z���kw����v�!�?�o-��E��>e)J"�$>�z�����p��S�込�Д7�PͱT(�q'�����Ϗ�)�QPc��OE��L���W��k
���2�E��kG?�`����mw�\��ߙ��B(�54�̾a��9�,����w����#��P��V�4&2���ہ5#;�5�P�\��뚪a�=Z\�*�Y��/F����N�q������HB�>^Ǫh�Z�8mˌ�oH���nd�3]�!p�s
��X���
�YJ3�t�l��H#.�a��:. �fV([��b��Y.��Z�ꌫ͓�f�����w{|�|��6L�0(i�h6ߤM"�u8N����U�ܻ%}�]�ˮ��E��¾񋋊}��	eu�;��5���p��
 -4��H�(�1++����.0��|���s����%�*`my<ʚ�oH�\-�M�t���?��j�˹��N�Y����	�7 �����D%=���kZ��gب��S��_��2)W�������8p�~GP k�"jMH�!�H;���(��\�̩lge0�*���q�hWm�tCՠ�wpl�v��i�<����"��翻�\��
G��RL���a<������S��ϗ������a�ǫp�
st�; E�p;W]<�;��g�P���Z��?�*��s��-F�y��S�̝�_���=g�䧿b[mb��U�-p3�=�YS���G��%�V�p�(TOn):)���>��h�	��g���җ&���P�B�6���+���&C������u�|�v�=MKCA[���q9VŒ�B$Q=���y8�n��f�u4�~`�[sd>���Lsr�b@Y5�0��O�b��-�c�0c�1D8t�'�٣����?>>�����4�~2-kR�l�P�p&�6�`8+ڧ�5A�~�7���yϩ]@`���C���,(�:�eə��c뢧{׵eQ��@ɧ	� �1	�h���rn#-��b?����<��(+��G��J)W�_�:7��:��'�QO�����*Zߍ���O�l���]����'i1+4����Mo  �3<�6�V&	̏�VV"�K%9�}�-)�F[�>���̕�����ۙ,~���E�j�5w6F��]k��/}
���^chsñϨ�DOBM�H�G\���EZ٘�2�N�J�;OF��w����$�u+J��mS�Y�@�O� ���+2GJ�6̓����w��7܍)�X5���dI�,s���	�$9�2�j����(�v��v�8�6&#��Pn�0:�F�Үq,�8
d��Ӏ�X(D�O	�I�]����= ��0Բ�%���JKC�t�v��ܢe�J�<3�u+�q��y�i�F?��AE����lT�_�"�DF�7�J���y�4L��p�jI�L� �p'm��* i�kT&l˥)~�!f��xXK�&ܚ��]q�ih�I�#�@����#��f$�X��Yܐm�W�2w�| v���O�?];�m<�'˱���fg\�Y"�_���O��7��|�z��WB�h���ח��h���\i~p3r�-���9*������t�0�sq�؎j�;
x��|<J]���}�|���4XhT���^��u}�$�Q�n�P��c��a>tbv�y/L��$���'A"�SH<X��G2�X�(P\���	���?�㦥)�Q�G������*��a�JSHVkV�f� �Ϗ���ҡsI�Q�0�t�D=^�-B���e�.�sr��:,��!{�se,H)Ot��YT��"��S�cO�pP\ͽ.pT��<��R�:W4j"(��W������ ��\�C��X/��hS���#C�U����w��C{z�!�3�/_�*]��0����{�$�N����fg0$G��4�r�N�O`/��[/���QRp�R�Z�ʶS]��!�@#�+cl�X�E]l��u��-I?����(���^3C;:V����k�'_?�w��N5:L��Ѽ`-?gC�u.����y}ü�����ﺚ��7�!��(�*��P��v@%x��A�e��MW&��6:�h����l{(F9�k��f5�=m�J<����Kʩc�[/�$
,U+��2�k��D�T_һ��ˋ�E��N3|?�U�N>�7i�?�w�לc	k���z�tT<�QX04�v�''*��B:���R�,����`��NK�5U觐�B�@�Q�D6̤�"퍠~ �*�z�T3�5/f����8r�l�B�R51Ǫ���YA 7��|}W^�8�}<<�����z���g/�]y�7vx9oXl�<��t����4�����\7����{���ܔbk��/�wSx#@1�i �x�J6Rh.X�/�'-�'6��9�&f�@>���'���
+3��{�s�3�L:.����<}^/��+�	�n/Z�N'��7;��6	�3���cz���Ƨ�9!�(٥O6d�D3n��R�d�!#!?��^bo&��ԛ=�;A�ݲ6��$��~AR2-��[��rhI��
'��~P����V�ŭ�}�h��;�s0��@��[îkFe��T~�U��"�(�����B\�ٳJ4)Y'-�^SɅ��w�_��E�n1��iV�O/�\��Ҟw/�JuCg)s���)K�"%��h4�1�_�z�Z��r'���D��k`�cxqb&�c0�T�
��H�G��k�����[��v�{�6^i)�ǐ�{��e������73��G���mY�G�����iqy�1�n��B�
�}�y��tb9��
gth+g��gU�kA�ŋ� 	Y>Ƨc�go�l��7K�f��h��J�i�PozG�H6e;���>
���At�p���!��9�%��z�" �K63�On�ke�����'4�Ĥ�b�]�4�7���SXw�*|��Vwdh�ڗw�}��+�LZ��+ҷ�0����0v�J ���!���m|'��(V����'�dx�L	ƴ_�>�B3�ffZ���"�XW9b�z-�-���K�NfzQ��o��t�J{#ν��-�g��9�/ �����d:%�'��c,���N�aY�[m��t�;�e�i�8�p��A� A	��I��,ڨ'	�}��h������#���ɇ����	|G.�0���'C�{q��MR|=�࠲n��V��9�6/&���E-%� ��|A�-06�4��7�8dK�B����(p�3�� �2TKD1�#*������e��s�H���p�ˉo��Tk�J���~f��aw�Ss�����;Q[Q� ]ݏ',�&�v��A���ށ��¾B��c'���:�=ԁ�
<�Al��)����򫣱���|g�$&N��ǵϿ�6�A���Ʀ��N�7��41U�MFx��T���+k�Ty_~ķ�0��l9دRb�)�SO��Fp�94|�Z��7��mZo�X���7��}�<$%�N����_�p�m��.d��d?^b��'� �)%�����"w����z'���}�����qe�a��F���s���ҥ�!�%�]��O���w��t��8���Q���;T��X�����jJ,���Y��o�*0�Y�W	�9Ws�\��oQ��/ZH��F�p��LN���Ž��%�cQ��vB��ͣhޫ��ދ�1�>{�&��3K�����@È�DS�j�鍲���m�KO�1]�n#�Ц���N��, �@��X��9��৖q��\���C;�nc���6��^T�����T���@٘����� y����˷7F�Yʒ�ͅ��T��Cu�־�����.zͼ,�H��Y��i;o.#�	y�$�����'��%���^*?������)xl[qi��m�rc����p��t?nE2�W��p�&��˚��G��"�G���FB9�>[��� ſ���td�|�/��V:_�f;��c<3�׍�BN�loQY_K-������.}�|�b�)�;�	���:�˗��k�X*�(�J�ŋ�)������L4^&"�⹴>�u����]y| �����Se+i>��R`;֙K�==uP����2Z�&e���X-�*&�cF���e��m���!��?�wtMa��f��:"ǽ���7���M!e{������k�K�^�����jt�7�.-�N��@b�ϕ �ۅ�2��� <Q�m�Ew7V��9�Ŷp��д.�A+��:��ĉ��Ԗ�wr�k�sj��/�Dy|>��|?������ ��^��W�~c���E="��h!Y�*���@BB�au��.�0������*�����A��GF�"O��0O#h˧����	����	ߠ�oY9r�Z�X�I�!��H3#�9<�):�e��"��&���N�O�?�w�
�rx�Ϝu�'��2�-h�І���#��q'`C��g	�7⿛4`�h��Ă�i��� ����w���zg��Մ�l{��Ga����b"Pꮏ�:d�q B;:��['k�0��"{}?���(_�iL�"N����T�F���ȕ_�&a����::>��wJ��Ӭ��X�����+p�٘�b爤��T6����v%�q�����*�(�����⟇���)���{F��aΒ<z����O����5��À��L�-o����;���Z�1%�f�	����2��Nے�Z
D�_`�/�_�";_LO}�}O}�e�����/T��V��	��͑m��<�IH֠���Y��yi�@���@���,���d�\6`�<��&#{o	t��Ꜿ�T�̏�)����b�}}�]�)� ��n�:(�����[۷%/��"/��Z�l��ł���D;㜕`���N�c���,���7�GB���%>��f�D
n�~<�ꠕz䟓n���9H�!��[���ʂ�c���IEHů�7�Q蜴P����_gc�ukQ؝}��AMm���3s2y�8��e���2�����;Q��͍-D�`�sO/b��9 mӭ�����b�
�-�+�tS<��|\L������d���i���/}z�s��P��A���G]�t�.>0I(���#?���ح��wo^�zlO��):o��ƺ�3�ص�]O��,5�����<�$��m3��9�x��'�d#��;���ZOY�����@���H��;���3d�u�d���?׸.|_L�[�&�j�`�]��3ؼ��/H�ҷ��R][6W��Cc�@�vb�(Fw�'���>���9��4-����ߑ�?��P�D����/ڛ��d&�9 �	э�twz)쬬L	i=mi�����5�_	�v�����y�s3���yz�j�w\��������y�6�`����>�D���I�F0��u�D,4���G��d��f��Yb��y@��b��wVSJ�ʂXC_!<[~�_�=FQ�c��o��î�7G)���!��I��V��v�������~C��Q������,���Db��y�%� �� �"����#�O����R7|�w8�W�>_���:ЈU����M3"�]>n1�J�sߋ�ʂ����v6�٥����9�%|bX=D�������<�v���h�l[eVs��a�#!	��_ �s �˻N�@�U=~*t���ğm��X�H�-�{\�4��-o	��b�d�E�n��Qk�����ӭ���**�Z������ñ�5;�Y-��O�A��;���)�~s��o��vg WD���E�����y���N�"&<(��-t3S�ˉ���$��0[aDn�qp;��f���3��7��Ք�(�i��sx.��V�4�M��;�F]�5+�[m(͕A�������x@�$�P��YP���
��t�6�z�E�38�[��e��gR:-c���ˆ�,��'3:Ix��8�����O���J;��r�&��8�1�	��D<<{]mڈ�`����2K�������2��P�3P��@��N��\_(4䤽U�:�~�adi�Q	�Q��:"�S薉�"ڹ~�2yw����`���(�O|�c *d�RK˰��sn}��	fnK[�� q45Uj�7�7��ܱ��1⽈��4��ε�s�����[GJ/�x�ퟪ4����]C{��k���ė����K�A��Zx얼��9�b��=��R=���X�����6;�윭9?��wߥR,F�ϑK��c��g�5���ڻ��UE���8�g	(�������F�(��X~|2�&�n��R��ے^���f��f��Hz�t�t����hE���󿳆���֩���y�&++xa��a��!�_�aYw(���X��O���+R�Lm���kR�n��2�O� ��|`"���|�	�u�Ċ�GGߕ6gc�mgUA���Ѫ��f{��V���P���pPLb(�q�<�z�Y��O����ɨ�����f�ZL��a�P��,�ʃS��Uh	��=���j/g���o���X�+��#yH]iRz���&|�H��Wi��)j(�������U�'*͌��ğ��l�B}�u��d޼y�i��)�G[ ���{5��Gt�60ʧ���㸘MT�b�K_}#Q�C����0��7���3i.k���O����
��r���� a�>g��P'�n���y�!�_O�dh* ��R� @S���`���!H���46����N��؈�Z!|4�0��l�I�f�PX4_�ͥ7�-3��v�:^�bp�k��[t�U�����9uTf��� �Q�VDV�$�$����ձ���D��]��S����bf[��|����]AAje����؄����!��V,�M��o�TdB�&����N��G�0�k����D���/3��A�!�6�;M��c:��߆v��q)���_�@��$�1K�]� 
o�����4��^F�f�7ac ���y�~�ኈ�����U��<���q~��I?qu� ҅�|���#"�9�ٓʡX�38�T���ѵ��d�������l��2uY�υC( 5� �7��0D�}a��PA�FI�>s�&I�R�g��/̜[������wY��qiF�#����L����b��|��+�_�$�Ik�D������e�����sU�k��O!�����U�M��F�� �n�ԟQ�(�:���藇���:�)��zcRJ�TO�OM���X����ho�Yx�O�ķԢ�|s(���`����1��c`����E����'Y]z�::^�&%Q��3�ܓk��VUGM�X�Ja��y��'j�f?�a�n�0	J
*�D���S�+����j~�7�;߀
-�s�Z�E,����������}i`�oD���j����nkSl�A^��xl��,���`�V,%&�<�'�)��V_U����v��0d8������-�c_�O�qL2�z2|�y�[�U����g���  ��8��5Џn�ܐ���_Io�D
 �a�)b֚�Ra4��^I*��&�=�ͽ�|�7a�4`�����&,|�K��-�?��k��ƪ[У�U��6Nŵ���T�V��d.j��M��v,&��m��)��u&�p��TnwgP,Ӑ=����YqL
}QA�bd$Aڦ�,=1|�_���+�)�s������j�|a�ǘXM��1���n�������~`���b�[}������yU�}H$�����,�Hm������חyKؿ Y����Z<Ã8
��W�G���2q�� ��$�S��zg�,Z�6���i�!���r�����/���Q1����x�D,��ِ��ɶ��O�޹	�� "���oVAc�.�P�1�z�ʏfrYiyt�e #��s(��������4��Vi�0hO޾���%h_aRWDR�����n"��ȥ�5^��6;W��G��5y�۝����(.�GCKPI7�s�<����麺��۝���e(q>�ز��0�ϓ3�H�u�Dr1�I5��u��R;�!9;�x��_^<�x¾~f�[
�[g�~x�-��F��r\�.����##�,OK���-�^��s������@]���W/T�T��HmaY  =�4��>��duڮ\Wq����y�>��8�g4)3}��2�D&��^H�֢k,N�7l�o6|��Y[�^*/�z���4�$�Ǽ��X�q�3���tef����)��1}�3�D����3��_�]b�Ù��%�[�QYٛIG����D��N���
+p覈�+HP�*RG����P��<�G8�����o�TO5^q��m��x|��Ĳ�?E��FX��a�ڦ���O�w~]�8L���l���O�����X@�X�Ε���LKkf�fg�
2'�2�K{�-�Tyz���G9	w�),T���_�H^C�uw���|pJ[�����kܲߌ�����3s��y�����(�RC-2M�aD����-�Y$~���!#��������/D�0����a� ��^�"�4�J��Ȟ�r���}r8��[T^{)#4�W:wj�������7�
�Օ`�8�:�yS�W��?�W�������K 9��Nn�4 �}���?m����4g�*�D�V�+�/��K���'C�v5
p>�*N� ���A������L֘�WZ{�[A��?.u�,8I����ˠ~��(u*�u��c��#��V����^7q�%W)���s��h֓�-�#5^W�����lJ�j�m9SQ�pl�ڿ_�D�=h�?jC�)�:��i}�2X����V�G�a�̭.`�*/<��Y�z���j���x����>&h�3�b�����a��C5$��;r�k�\�i�1�w�����0�%Xp�a=�҄��\�@f0��R�X�?s�Q��0�Y�J�������Wd
\�!yM��38�Btq��,��l���~������~.e]��F?:�oJ�� �d5v ����0%��w
	�,e�[\$�LISSl|;�7�%x�NY���'W�I�z��w�f����5]A���x�H�C����^Y�m�6�W���]7�V���<�5Q����8�S����[C�D+�:��s�'a	7�"|�pR��XD����j��	Wae�l���b'�y������2���P�cdI�1�P�8��vF�-���| �-)5fc#{+�z-6�����WZ�E���۷�����o�E�p��~��Ǥ�݃IW��G��\��w��,|�ʽy�2��k������g�W�9��6w`�7��_u�����ɰ���R�<0=#O;��g�
K�9o���n`X��z������7I�tY̟�����~�V�k��m4$���%��?�X@,��$�=
�L�$�54���,�(���~��E�	��[A���$�S;Ԇ�b��w�����3���TT�*�mrD���(}�!.�2����K��S�i0�]�>����YHp���)W_�ڇ��N(�Y���l�c�.��U�M;?�:֌{�#��ĳ �:[�L��M"�6f� �ף�"lͫ�^����0�7N������f��-W�\�=���ʚ���o�U]�ǉ�7�$��2��̪�o�M��D���v�
!�����_�Nˍʈ�����o�X>�~�{��	�)W�%�N+�[{icL�����5��7�1��R��C/d��q�,�(��z���W�M���Bq���S4�|N��;sh
Ì��9��r��֎o��F�|D����fŞ�Q��=
s��D{r6�T�z�,4Yz�'Yԡae �b���z��phO�H��+}�E�%��2L���O`'�L�`����/ñO#�)z}08-'��NH�.�S����u/��G��d>�.�$�s��ٲ}.*j�??�(�Y�J��C�έ���f
JR}��-"k�	z�U��gT�z�g|���/q�/QF"2�A�
��I
(77���ʮ�8�x���7%�Q$�xe-���I�����l����.LIX���mj"�Yíz8>�A�<�qP��$���[��Z>x��왂m=[/�lCe�"��km��o���$-�x��#4E#�ڔt��<i<2c��}o�%�I����t�2u*3�l�Qp4���1����P��C�Q��;�����7�=
N �����KGg9o]��b�c{��W�2�ա޴�����(K{0ˌ��a�S��W��7�Ey��(j|��12��I6�����:�'���n|��S��O���/��T	f2O�8wn�$�O���##�KQ��pX�I(���f�	L̖��ja�t>H���pR��E�(vb��㹰�\D*��KL��D���G'F�1.<�L��I�#�ڛ����.�WQ��a��y׏n��fz�Q����Ĕ�r��j��I��󦜜	���
 ����WA`�IH�_S���ҎiVnjo��/`��~��*&Z�G�Oif�ޑ����Y�����mUQ�c<�[��B3 [K�S���,4K��1��8"�>E?�9�pebv���X@n��Op,��7�'����!l�'4Bs�L��J$��nE�(�����N��oK�M��a��W�Ā�KE����.��H�f�pA¬L*�v�I�}xЕ<
AK�p�_cw����ɸ��\�4��M��a�������)׵K?�Ʌ�gU��FĽ���LQ��no{���ܽ���W��U��ʔ�^��XNt����'O�N�
咪���Y4�^/p�~��f20�f����v+-�X���&w�A�"	)�10�eF0K�n��%z�sL���E�K��T<6�ehb)��?��*��T9�>�����:�n��?��;5���� ���HB��,�Ѧ��\����dwUW⧻d�0pZ���J���0��{���G4p�ٶ5zz�kY	�tԣ�1*��x��<c�^������ģkW�1#-_�D/��OUP�Oܒ�[�6	، >���li��f(�<�RM(2�b;����J����ny�Y�G�.��ib�H�2����j�2<�)L_k_�F��m�]bN����=,��{�:��1�:[SQ�.i�����>%_��SA�m�v�8+�2��[���U�\���g���Er�~�����d���`�[E�Ri��Է.D�eVV�%��W�O].�E�>�c�9!�K�Ѷ�ӂj��H�ɰ�ǎ��O��l���5����u���ad�ϒv�w)P�?�T����u��f<��y�D_-�;NEI)9#��j����}���x��EK��͕�;��!��t���_O���l���X�����/��2�I6��W177�����C��?}�U��.؏8v*������_�"��8���>~�n�c��`���ٙ�]��	����`>��?ED��D��x�=���T�;+vDS���D�r�Lv�ƍ*�n!�rCTQ�M2-\��.���Pmeһ�xv�p#��N���X�#֘�?w��C��sLz�9O�n�Τ�17��c5(4H~mςr/m��us/GA}�K"�'2��Y����C<�T�oV��V��s힡%��x��!��;��DЕ\~��Pέ�DC���2�!+Z�Fk����$P�X�A�#�r8��[��A��+��Ě6�^�2����8�JM�- -�=H�
xvf�H��Sèֿ/�$_����΀*[D��+��E^����ypP���p� ;M)3�l�����>��b���� T�ad6x��B/��;Od�����|��x��zg�H[\��TU?zm�;���<�`�}s���܊c�����ʾ��H�y_�g�yItZe���c�%��:�X�Q��Q�d��6����]=�[U�峭����{�V�+[�b��"[����SY�3��ӧ������W�����P� ��|��12w�_<�Z5�ݦ��*���S��R�5����G���ݭ;"�1��]e���t�g�
�Y]&���Tu��MX jE��G(�]��C�����59s�_�IE��wQ ��F���9H��ɜ��~�sU��oҨ�\l!�lɥ&�_[�� YI�WGǶ� `D��f.��<YS
��#���&8_j�Hq��S��,�W���^�F�!�� ��J�����2�'�2C:Ǔ�(�i^X���
a��&����e2#��"']t�%��@Do�=������t����rs:����#�K�]/��\�O�Л���Z��.4^A���珿ȥb�9�,xvq�\� �ןx^Cw�Ia�ukħ��J��xD�	[v��FuH۪�vtؘc��RQd��u��U�z��UԵHG4r���Y�z�u�����ᇧ�l��RO/!1��!����ђU�Ͳ�4�_����:�1v� ���bk�#�,�C-3���\��	��j-�T��ӻ]�'�M��v֊׀�_�B�����*�й��~%��u��+[�Ꮀa��;~??/�(�@��� �H2B�+ǟ�7�rH�J���:ԯ��%'���^�]o�	V[�74[���;�(N9������o3'��RƻM�FJh�5�ҍ��B��p:��#�\�0����9V��2®"Qy��8w�x�bk������%�׉"�6Jt�=�F*NUwT*P��1.��d�ֳ�^S���፤����Q��TPɽ6��KY��a�gΗg}���t��T�F)W�qX���&8sE�"^�����w���mE �zE�ϣ�`��|�/�s�ݐj;�Cd�R�[y[B�QV�>���&�7��ii5����C̡���u�.��N#�ѩ���j���Y�|��JxIoE��߬���.(<t��n�P��kB�mu���_���������J��c��?08*~5v����
�ƭ��*���Z�_�k�pv���^�+�G�v��v�~^!�?�/N�o��7̂`�}�� ]W�5Ftԧ��Z]:G7p���r^U����*��� ���Ѐz^Խ����������7�OT<�3|H�a��G�������ӓ�~e����4]}	̵ܑ����n� �&ì�����ō%q	�S�ƊP>N���UG"�u�M*�ۿ� �t����O��g�ء4B����2�P��=�Z�^3q�|�.b*oq�c9o�j"�7AOw��̴Q�F�w�����$g��48�b�jUZMd,������m���PQ�O_	O�v`ڀ��v+w�w�2�OL��R��)[�`�Jr���v	
�~�k4�Ѧ��5?�r��s��H�`Dio�n<�!�����p+��_�h~Ѯ#~j�C�Ub�f���E���ֽ�����k����>�'�����R���c 
hd��A4rF��H1���/��YT�/�Յ[{���fF兘*ZQ��75�-a�������Ո0?��_��
�UM�@�2�m�qV���4��0+����j��v��%Oe��uE���\�D^9<���xh��^����rS���&����Uo�k���K=��B�
�#��L���aЕ��7����@"�`F(ï ���Hȴ>���Y�s$i�������y��0������N�W��R����->�mӃw�/�x�ǆ3u����}����`~.��i��J�FTȒ!�F�Ay��͍���ʹ8/����*��$}*����BA�:m'�̖_@s����C��kg�~��얗>R��;Y��]��\	���
^E��Ϋ��Qj����|P��s&[viA��5A��okk�dT(�7LCA�z��Z�2����
>��cgfy�d��VR������P���.?},�b�&&N��9�sw�d�ƾ�����P�&N�����zn�#�#��0�+̩�δ[�5���0�X��sj�6���Ҿ�Ejkt�o����� )Pd�Q��A�o���#�#n�
�SUV��.�R����S����>K��0�C�^���+�r3J�E�h����&P�rߗ��:4�O�������>#_�y��;�j{������-��̧�WC%�O{e�B��������)b���[8��B������y���iE�2P�Ŵ��"��K��E��1Z��`�2���᚝�ù�kN��7�+*寕��`\�+H��*5F׎�'"�Ұ�9L�2N�;KׯU�{w�H������xd���h���"�]j��,�s_�Q�9�Rͭ���7�	l�]q�ҳd�w8,D�Le��֯e��y����Y����_u-��*'��3̒�����_�@�?G1����Ϸo�[�)g�"����4_f�x-jO)gK��\*Ƿ�9"S��X��������}{�Ȉ����фt��(Bv��@iIl���9e$)�U9i`� ^b�H�딀8���o��Γ��L���߇�\�d�SZ�[Q�O�ua�j���7��5NqU�����W3���=�L"/;��'���A;�|5Op���>aC�ɽ\��;%n~�ĸ��A#�M�1��鉋٧*b3���U�3��
z{����W�ݐšN� � �Q����t�W]U&�Y�6u1c�������n<��K�T4�Y���,<�����X�O���n�^��������c�<���j-� ���3���H"���;ej�BQ�(�`�}9�*�J��f�u:�oMAQ��NMk��g�+%�A77���SE	h���]�d�p9#ޯS�M�]��6��z7��v��u�s�Z���m��`�:���q�u8 ?a	�ĥBfK�8d�E����tն#�+fTf�ޯ�#�������&߯��4(�"%݈�4�t��!]2G+��� ݥ��-�AA`����X�_����s����\�:wl6���gf�� ���w��`���^���B�)� �t��q�L�w�B��A:�+	�MX�,�?�
�-�J�X�E2��ɽ;klV͇.�Ҷ���!�p�P����L�������� "	���O`��ȿs��40D^���������¿�Z�H�d��:1�@���x';F��.�أ���f3����U�3�|�q�7t���n^e��ݺ����3[�E�+?��oL::��"]��po|uW����ފ�g�����F��LG"�Oj�Ҁ�ƶ��Q�<��'��ճ��'ܰ}���������8%��r
x	�1Ti����H�<�l%�4��Ǧ+�pvd��wh�EW~~v��,��
?��W�ܭ?���O���w }=p��m��v.��O�����%m�n4At%χ�wi11B�����ޚ"%v=��K�1�`%ھ|�n��-YO��G���\�^�#��y���ڳ)e��}�"̿��/7���}��t�׍�P�U�"+=��s%+2�=9_��\�?ɔ��2�]nئt�mJR� ����[9+#��06G� -	O����i5�7\��jHD�L�WO�2./�^�쉔i�v��K��N�!��?��m��6 �=�����0oKQ`��C�&_��_��|3h��֬��'4�����[���PXV��P<A���0U�M�plλ�9+�؛�[(��S����iW�������<(
�T%+<�A���׌��Aɝ�;��+� �7�@C{�#)���|Z&�����U�H�fNnZ��fb�~2�u�'��T�����eJ��toW�zH[�Ro�3�Y5�3�+�mqu`b	���o&At���e��N��l%hS��^�?���B������E&�`$'�����2Ա��w_�o���׾V+1���?yD4aW���E����2��N븙��:Nk�)�}u���,~E�Fs&���[����ͪ�ꅰ��6��`}����K� J*Bz� �$&�eAY��e���κ�2f�Y�/ߓ�j�PP���LX��t�+{�)�x��n��E��
_}�� ��:r&g�
N?������Y�� ]b��~ TI�g�_�WH-�S�>�Mm�U�:)��:�e�'L&?Bł��~A�#wV5�t�I�@/�RW��?��1�e�GP�&,�LS���Ղ�Y��~+^�0�����5߃���>�o��o��E�����W���û2�ʔ�lYz5����?}����%��Ǳ{;��?nܗkѡB'�3. z�B�Es�%�'���������~�R:A�J ���X¯�T>�V�ǻ)�����s��_A�O��I��/��4
\���N_�Nɔ�
s:>��_�睍��p��R�����P��o��m��L��WO�@E@�����e����.z��/@�/=�]���Y�좇�0�Ue��i�B�zs��0]��.|x�G~Gԁ�¹#Kb�G�#/O���P���>0io8Eww޽��hg3q��$����1��w?A�_��%!< �j���v�5����fs�?^�rͩ��:����gD�ޡ׾dX|	�%A������P�uࣆ���a�BE���wD�z~�K�g抨�Yc9�.���-���%�[%��_�I*R�c{�{hԝ���Ԝ�!π
�qw�?�S�����$��E�?{<^�����~[�\�Qx&���-�n�MV��Z���D���_ ��ւq����0|���8�	��t��s<�����7^��2�q�*aB4��~�?>��������:�-�-�u�)�<ﲽ ��QE~c�n��Sz'Y2�XK�xPWB��� n��!R-ǳ�p�xb��I7�v�t
����'�F�dt��?t
�Ջ�#��Z�ԍ�8�%�9���^����^�J��/��~t���r���@��b��݌~���7�\�;����9����=�q���.�����i'�8%�T��Z�x�lrg��s��tÊ�Kh�G�r�$���'��77�C�:]��~s�W\X��?6кo�_��)=���6zh���?�}���#ߕ]�v��S\��ᱯt)��+� ��r/����iOҵ}/�F�i� �+��h`����l9�l���P����xn,ŝ�o�	�H��F�d	��6����!�U	Պͮ�+�Ҹy5r3V������./
K�g:�ǜ�?f�߹-+� R��4�a�s��rp���+q�P[x���>>r�%�j��q�P"�x�V@`��.��;]��I�P�9xM�����S����	4~��}dT �u�9~�������bo���.���GbM��Hvߺ��2���JLd3]�H���c��R� Y�$����N�UY�<So��΄E�n]��*w_&h�*�Ȱb�qr�&(�)V�n	s 3:�Z�_s��!�˙S9�l9��u�������qDo痄e�W��d���z��ˁ��8��i�B`p@I?ӂ��j�<I������U��X����5�d�k݇	���_	~�K٨�Rx����fD� �o4+�x%Qo���"9xˊ��~U���8]��>��}��~4/wǔV?n��#b�E�7�l�x�#�e(PFQ�o�����[�����k���+�yH�R����poP^�C;�3&��1�ZU��.��|/��?bΠn_0��Ztճ��W��z�ԿŠ�FYʜh̽�^�4�WD��Y���'��کW �ѝ�A�W:oVUC��� \�/�g}p�":�!I?�rs�VY(�H>�}�&��D5�Ͱ±�ڿ&<��⽩Z��E�˦�G���/	#O�~�*��뭅�������L��J�U[�(1L��Y?MW�I��~�MM��nA��ȣ��{5b��4��!�#��A��/�B��^����C���^��%���)W���R�q��c��WN|��Ak�6ڔ]��W�~�*5��BQ��C/��eQz�@�1sm�O �ɏ{,���H�K�_�lc*ƃ�/��'tN��`�SL���"�ѱ�����ҫP8���:�q@v��A��z����Ĭ�+Q�*RJ�%�����_�c>�Q�V�߸�᢮n�D�Έ+_}*�, ��@������[��F�OR���I?��x<�M*h�	}�2,X��P�3�؟��,��p~�$r��@`.F���&�y?�(��3TA̰��{�xZ�t#���Tʬ/C�#��R��7=��g|ů���BB��	'�$�?�.��X��j�^�\��1]�y�g�Ŀ�j ��6��-��
��c�\}��MM�R�2����EA�����l~ۆ���K�xC��5=|�k��N�$���+�=�
��vY m���D���o��:bS͌���o�����{v^�\2�����MMQGx��m?+�<\�d)M9�m� >�z���&A��;�:�	��|$u�F������Ԡ�g�P`뢉��IsǼR����O8n�xi�7��y^����3G��o�|��f��(!1�U�߳eWS��*~q҃�x��Rʄ@�L ��U��?�Z���Fe��?�p���?^�|'�ƻ�:Z�ʏ�~���N|��i��
��a������~ɇc-r�Z��-��r+	6��o���?EQ�6����]��]���OmSD��h����!�Ԝu�(���1����v�^�M����:F��\�O"Fq~�i�	�D֗����gW^쥚a����g���)��������&���9�"$&V��N`��e(��T[)��Vpoo�٫��I����z�L�*��0�}8�=��p��Щ�H=�Ӂ�숐,4��gx����ie����Lmo�a�Oĭ�9��͒D�<l�,d�UPNëm�'v�;��, 씰 o�?{�K�͕�?'���y����=/������A�@_���5H�5�P����W�׀7�?u�a�3e�cf>԰�ܮ:)��?��`Q.�J�`;
��D�z��z�Ļ2G�e��rk�!�w����{��S�8���	R��´�&�,�T��`N�ı��lp�NI�!jů��P7I�od������\���T�ٳ���þ�� BhpO8�GQO�Sy��9��ÝR\��Ǚ���Q<�B-���(5�9L�cpXs�Ƥ,b^�y�H�*7���I����d��}�c��Z68��3�E���X����K^�X�|2��Pp"��qi���e$��=�	��݃��z���<��b8����CƵ�S�(љf�bSZGmA��@ �"���Daqa�j�kP�Ş���R���|�sQ�f�$(F�Ͼ�G^�j;�S�To��)�L,��b�8ˑ�\���%[�qz��#�Ku�sAo��`�m�v4p����0y�cn��`�s9�{�I��C3�q	�����S�����s[�%
F�������h�_��#=�;��]�ZڗI�DOٖ3O���3.��y܋�GǷΔD�D��o&j��,�Rt8	����0^�]`����)X�N���R���%�|R�F��Ԓ3�y<�2�/��?��d%2I��~�W3O��t����T�%np��աW�~;w�!<�M��R%��`�y���G�PU�$I �@~�DA��w�D�,#2�J�}�S�Ϲ��gWs�;.X�/(���_�"ç_��lދz/��M�µ8�_c辖�w�ܜ���=W��/ls	9zFƽA���N��V�ҝ�g��5�:)O����,e�}o�$H�k��AS3�����m"]Qw��+��n�����%�z��:0�w3�z���FdX+�}���d墙?���ad�=�%1%~NF�<Z6�]���s�z�jAEtf��+ys���o;VD��U��3_3" ����V/��+ŧ����̵�Qi�2|"���P�[�+ۉ�dҚ�Q�h�D�����ϑ�a��|��O���J̯^�K�q��|��ּA<+GS����YQ�f��D��h����� �Q7��<դ~���r�x���I�e���rԲ���x;��-���� �i�{����7#u�F-�}��w���7#"��]���7��޵�R���h�F�1������l4����?�>�����w2oR>o�r8�v݀L���u��yҍ��4�M �'[-����%�*x,p�Hٮ��ә:��ý�ї�g���1�J�d���,�~��(�Ga�8^N�%GkZes�Ǿ�I���a�!��7���oܾ.��u<?6xE����ˆ��g5��~��L8��XT]MyK�]�"݊(�Pׇ���4��h��v"�ػ��Q��u?��b��k>B�[97%��-ag,
vz������t����;�qad
�\��M2�5��M�pT�nآ�v����R`�;>u�6���(�u��G���x�o���!bX��oe��U!�gdl��<�]l\OI|��>��/WG��=�'�YHVK�q��x���8V�+�;��@�l��M���u�p��A�����F�9�Ä^�(�Z�M�Y������b[���:�w/�}A��a�Ӱ�o�$9�ż���u��Tlmf"�� ��S����ἧG}�6��0<&~�lFݏ�wmU]�I�u��S�%Nmr�4̉�@�8�Y���Y��!���2���NI��&����06�r�o�����:�V���B�J�|�w���I���V��b���_�p����}�|�h%�3-T�?1���W����a��+w��PC�D����{NO=���)��/[:o'���g�X�#�3��A!�|����ڊ̿��|U�ƻl:�RV8U��[���m�(���8�I�U���5�D���@I:�)ڏ��x�06��˘�Z���h�ϯ����Zn�����Q1F�q�u���M�׈S�[�k�u����)p�@�>���������XS�j���9��L�`n獊dg��ɬyȌ�?U ���s��"�q�ս��l�ǅ5���T�7�{r�1�P���oFM5�����h���N�mN.&���ظ�7�jojm�i���H6����%ݷ�MJR���"��iE�O7��8@��1��6ק����56�6?�dM��6c�q���>�3�`.�0��0(r[�b"j%�f+��[2��Ŗ_�'�kB;b��P~�	{ǎe�#"4/�-��@u*����p�J��s�2� �S����D��CM/.��b�+��t9�02{LE/Z�ny~�	����ԡ_gU6����&���Z|tÛ�J��*�g�,�P�Ŷ�����ߞ��=����Z��)|w�2�0&o�>�Qc�sD\�|�ܼ�޻o� u��}��(��)�?8�_#�����]���u�@�ڝ��:��5��Y�s�@!�}S(��
�R�b����L �43s�<�(����ӥS�������Z~@�-�p3=,�2��/�
�Y�[��_�+�<�=��V��$D_��U�O��Cb���ݶ��"�4>ok�	��[�^�5�7�|�@�W�sXAR]V��V|V������"��\gԠ����9�'����E�f��Yb��Og��Wl����~lX����<i0�-(��\A�yݤ��d�,�s{�/�t )b���gP9�޷��K��*9 ��nt�s}L��}+-�24��K�ji���_>�%�ҍ�{�$l5���
-��.����$�E ��HW'[��i`����h�C�c�6dN���޾I�������t�'��ʱﾗ�
����|҂~�8
�y\*�K�Q^� 5��A�e�z5�����y�Q�Ã��7�,��������n�d�f^W�|r�5S���}>|�zoY~1J�'P s��9|��	�Ad��O�bu�Y�T���^�}��䄬7RN��F��	��h`{�<QY�~>�ƱF�!`�m�T�~մ���A�"� ۤnf���b�/���V���QT�:�Z_�*� /o�>�)gj$�� a��b���	��z�"�D[� +���UGDx�i��64��Z*���XE��n���O�ML5�ǂh2��9���@�}G����sS���t�0Ԣp-7��kS�.1F�W{���6�`��w���$�����f�G�9�<�0�B��4�?�,�ˉ�hM����f�ֆ�>������]1d�V;,��Ud_3�[������3�K����$���s����iI�U��\sZv)�+��'�gJl��v�����*?D�tF~�P�v�_����]�'G���v@[��2�~���|3�ͦ7���u5�h��4��<�o��Ǭ���9X:ӯ��>\�>�}?v�:�;� �V�A=-����*��,%�ah��8�}tvrAv��CS���x!�Ŕ���6�ċ�X<�`��Z�N�~���,����նY�Q�C��ؿ��ȣw:'�<�잩c��&O����y�{k��1w��	�d�58Ê?�g$�)�<�J�vrf�~��O��"
��Ks���ʹ6��۷�p�ȏa@p��ߞ�����Y����
���	��g�U����R�6�(��O>�/Sj�|��C��ÇAɩ/��h!0������T��Z��R�x_���{v?e���Dem�J�!V�d�|䡖@v\�����{M��U"�-w����!��ƭ��KYC>n�*9c���6��`���7���rǋ����_�y-�	��9?nq���f/�� �x�2��0���Sf97_4`A���TEy�mH7�?���9ߪ�Qz^ * ��aR�89>Wc,�D�y[�=M�7WQ�بm��X��!!.� ���`ے�6��l�L��8��S1E*�#���C��P{s#�V���S�����LML��\�qD��$�'"4�����4�^�����>Pb�n��n����@[���(p��@��T�-),T9�Ӯ��lM�� �Oo��B��/�~�{�Vp�W���<FO�/����b2��i_��s����Hk�	^�L
����"T�W�@�]=_��߈�>��_��C� �ЯE����o�S��x;v+��H7?�w����:P�RP��pΐ���P��%
k��rl��P�������xW3�F/�4�����g얄i4�5�n:;���'.�R�e�>Pu�ؓ�� �>T>',���o�E��CY�,�<H�,=w��7��I[�rf���8��Uy�/GMG�Mh��;��h�d�;ri|�S�6�����������9lð�9�����%�`�`��W5zR��E'g��BZ����#'��-�{�@�B���:�8��q\#/boC�Qve���A+w��l,Q�+�46mǫ�V�4����X Z��!-����d�n-|��~71�,�hUr��8oJB*[��Ё�+j7�<}2x����+�)�2���e�� �x!O��+��������sa����=��w�וV�^:eW�w�!r���V�m+�t'H����?�ţ,06�?!��<�|�~q��"=�/�br����`�Y���*�Y��F���#?vP��ʠ��6�8X|R����v�Ϭ�z�X�}E	���͕��E���|��՘��.������NfP/��)u�������Ƽ�;�� �uo	:�,�6����2���Q�!��̡:"B�:B�
��	�����X�'�'�p?�࣢�%���騻9����?�+ߤJ���^�j��?)Y���̒�GpGf,O�c,�aQ��,]��u�(k���D���~�+n��M��#
�k��0Y�����JDɥ��JB	:��y8C�^���x�}Ly�x�`z�W��nK.���
�6��"���<���J�����/��_H5l{E�W��������cH�IM$��|��D��Y L� l���	�f=�bd[r���)��WI=Bd�������b&��a�& �3-'I�9v\��a���j�C~K�u�/	�������'�wbA�y�ʽ��UP:7<y��W��$#��yGkA�� /H\��Ӻ��"B6.�w��V8bU���[D �����
����!����پ�M+��E���d	���]�/v[[��������]/9�v�CT�^��8iΖۧ��E������N��UB��+.�`� ؚܝ9��֘x�NN� �t�3�D΂ P7Gv1^��e�om���{'~����8�SP�e|b�=�M��Y�X|�)! j��t>j�����V٢���Ø������`������p�㺏�5��Eh��.]ڟK=����j�}ٹh�O51�@�h���v���ٖi����JF�z�w���=)�O�d����,?D�	@Y\�-k7U�u7B�*�ud���;??�:O�D�^ͽa=�<��^p#t�[ :�e��JN󯆬��Oz��o!r?��H�.�����EH*|���Y� ��`��ܾ{V�G.�����z��i�J9{�!�\qBt�lv�:
}L>S��.�O�p��`�c荑 �^��ΔDʿ��g����.�-��.a	�q�қRL?���Aȿ�/�}Vt��5��W�N��
<YyM��ɺ��g��d/2�7�s�E��T	�[ �D.&6����~GUj�le�����D��z��d���կ"������
�S����E��9�ߍ��iZP��Q>��ݶ64@ܳJ�mV�A[/č��mI�͜��9M��x�"��x����=b��^ie���+{�?��{A	���O��"#����+GE��{7�=�?��;���o�$6��]�h8�#;=ݟڥ�l8;
�<�#>B�S.vq4d�t^��r��w�>�&���`���U �@=&����uq%َ�"i �@�� WYE)�w;���Yw�$�p~�Re>w0o�X�+��7��� r�Z6`3���<�OfK
���`�$:c}(u��j�~�b^�'�vi��g��u�S#�)	����?�
��Yh���-��Ǫ���Y���Ӎ�u�ͩ�
����� H�g�J����d�:n�mJ��u��m�^�O�;�^ԟ�M��۾/�_�-� &���j��m��n���bچ�	���)u\����?��оS�(����
H@�1'J0�V	@���cGs��Gwi.�4���Z�ۙ��O]k�d	��TY@����*��?�p����`����!IOz��W�
��W�� �;c@, ��u�o*{�m߄m4��x�(�
|(A�\�0�䚊��/� j���{���F�,���������.K�F
R�|�b.]35��ŔTM�Y�5ju�l��=��=YA����߫�>�F6��@���d��O���{z��ZLq�*�D��Q`����g
��b�Ͳ����˴�d.�����jl������ަ�-ػ6f���{��Q"W:(��g�\0B~�n����cI",`�ͤ�$�36�m�� mys;;�;�t�����-i/S����7��Ͼd*z<�P�g���g۟,�d)�"X��[��Vf�%j����p*~�ǖ���]�yB��뾣�}dZw<y��Mm�`)/m�bd
݆�7��h�)���Q�~�?��W�p6�I�v��kJ1�K���ճ�s�����}�2�X$&��F����!Ӷ�"A�<^\;{���_��7�K{+=��=�~=U�/4���E�`@4����)��(	"�U�X�Z�L��m�7�nY�>OU N��l�v*����9�S�JL�����7[���750,�~�Y
���$H�|��z�dsb=���*�6_siJe6
�{���zj8���I'�OQ
O��K��-%3��oQ�3���5/����+�SM��
�����{�d좾��s�mԬz�BMvw��ʕ����i��{��6��[�n ���W���Ę��P _�e�I=xd����x�=��?0�)[�Ցw�~�v\��\'X.�2�7G��\�p"�PLhlߨ��L�)���9����wM:�n��<C���n���\��Zp��;��P�h�J��p-Hj��VY��������X9�ȗ�gJ.����z���e@��S7=�����	׋�2%�B�u�,�<��DzD� �,�ۦ�)�B�&���c��D�Yx�A�;},Y:�UINO�y�S��5����1d]��r�F*�ͺ.�<�&c�h��"��;�HL�:�W?�|ǡ��̚	��t>�H_wW�%ۛ����È�,N�O�T1�_���|�g[���
�^V�Lʩ�����sjw��%\����y�m�W�Dn�%��MyN;*�^���~̚$'�3H��xL&a�{ϬE`y�&���vk8|^�����ڏ��!Z}"��W>��r��̏�X�M��7��4�V$a̞�)����N~ɁxT�l��	mkw�H៳�����D���R�T,;9GY*6�ƑE�.po����\]n,�������A����|�AE�d�"݊y�� h0Q�<�(K�g�)S${7��u_4��w���� ���H��H��t�躞G�9���|��#~Xp%Fb)g�tgP��K.<X$!x�q��cS�|N�k���=^u.�Vg���z���r�.0%�����בŅ4�b�ɩ�]���m�B�*��]}����y#͋&�����a��P�����^�Gn��Rw�e ۽BQ{���+����t۬  �O�E�n������w��os�3�"����(f^k�|�kZ�����sD���^��u�1�����q�&G���
T���0��h�v��Txe(�;��ǾNՎA��dRO.oѾ��-HΡ�b�l��W�?��=.r�:qV�Ca��z�$��x��;�A�&)���1��!J�*}��������Maٔ���y�zIRh{Kc/Qn���3�����x�ܗ���3�}�$�ro5�\�0f2��xy9"���D�*& 6�O���K�<�2*i��8����:*��>W:���?�V��#P��"�ohU�|�1`fCv�a�<����ၑ� �� ̓y9\�&�/0�ѣ����x�_�U�d�3z0�<G
��xE�'_5|��椎��Z���X����"�>�������I��؟[�����[��9s�P�`s�SNo��b�Gv�C��Rԅ�Զt�[�HA��<�c�k$�3���1�vMl����.�-��+��'g�:���pCA����e	���2�J�_��	׸<�� �N���0�`��P	~�8	�y�R4;�=�VwL��j��|��t!:�3<Ʈ�M-x�|U�-l��Ax�~/r�T�d�:Wg� � Yje,]sߤ;
���i����W��S_�7@��O_����s�(7��j��es6��!�[$�;	�@��Z��aV�W��Ό?�'g�ݵ�i?Bѕ�6�E)XsKô�+��P��΢c��3v&WgKn�}@Sf
����#������#Gx�;��g;�k/7�� Z�����G��$���_qݵ|WA���7�f��'ĩ�o��O�I��W���DdW�?<�k�N�3a3�vhB\�ƒ�:A�k
�������W�{P{ʝ3)V�P��y�ܾ�Х�N��@�<hqP��Y�	?��LB	�kf�H��jc���L�H��9*���O�ׄ6��	/�\��Ö������cՍ/�R;r,�D�5<B|���J�I�a=�w�e�c�4B�~N��a@Ю�	E�ǩwLV��f��F��'R7��:m�����叩�X�s����%��_�;|~��{o�c��F9@Dr�=���#(��Y�=1���f�D*��n<"��D�[��V0�/��
��I��N�H����<N���sˬ`�S�b?r1��3ºe�;6�tk{�����u	����\���i���$�6�^�^��βBw"��ے �N�ک�R�^�:�]pP
������߂!�~�5m����EV��;��m&|zx���r��P\M۝V�D UR*�o�\{��Å�6���W��Ś� ��59e��(դ�84f��:dr�U��/t����iޖ�a��x�c������ld�[�
x	@02�F*S�E���3�gF��s�����9Y��ύ�V�k��T _��������vZzni�Oe��P~Q��m���V(�
����P�G_��~ }P��׹�(s��̚�dN^���k����N�A�ӗ�N��t�0��W�HM�%�}kI��YD����q�1�f�ǧn��{�gIrܟ�q=�n��t��3�=�l���*]>;�Vv]���J �*��m}gYlqZ�V�hɽ]�2�)��AĖ(�%S��b��nV�e��X��|�j[,!fd��Bwc�1H��V���Ϊ<�յ�Ly)s��I/R��UCE�=���d�m*�	�g���Q�6�T DSl���E�@��,y�U��:�y>�@�(��aiS��I]A�Sۖl!dh^��9�����8Q=��?��*Z�8�>���a~��Ob)�8t�[z����曆���Z$	_�Q�Ɵ{L$��1	�K���A��������]�GGs�uj5֞[�xuU<��_(%y$��|-����tez��o�,ҜIb���kώ�M�w�����f�Lg�-�ʿ4�V�0}?_�@�Q���
ٳG��S���Fy>��ء��<�"��K�����G��)����/�/\Dp��;l��7�Q/��Z� �I�+r�+��Lr��m�_g��C�a�h��<�7c�X'.VE)���6�jwS����|�_���C�'R�A�nT���1<[��/6�>���T���r�h����¸*.s�)B��:z����(����p�Q�9Qt�A�n-�$���c�����篤tt�z{������8����5�'d%��o�����GK	�ق��ٺ���7��O�m)��Y�uE��ތ�r�)��*�3���|��M�^��0�Cjv���������"�2����q�X+��"�9]q6�d�HiN�ZF)b��$n�t�� 4�}�c��G�n~�����&�?���^�I"�o�\>�U�E��)�t ���t���C�4e�Ȕ��� V�?�s��W_{e�U����6)��/�c�5*�	�<9&�J:����B�#�6&���(��=�\�V�,x��7j��c/��h��voX�]L>F�#�q�z��BLz"�1�ſ���m�	��Q\�Z0GC���j�����D��'.S.� ��CB *���qaHAٴ+��W�QO�4��l���U��W�Oc�O��|D߈��	t�jb���Qw��-]�V��Q/��+,���~�`�7�� �a�c�� s��}����^+�%=3ڞw�樷L+���y�V��_��1!|��;�a���O `�+d �|�B B�����҉�ק�0�*�|�T�B�H��z���� �;�*�4�@h�����4]����\�D|��v�h<_��n![M��v�Ut�!Q\{�}�6~�%�R��:J���k��A�r��Vc3O�����pƉ�(��@�ґ^@:�� ����$Ąx'�O��/w0�����{�dQ�GN>P�TW�W�\�\��8��
¹�;�� �~Tnϰ�r��E,@���6��8�
�b"?GM��pǦ��y�&��q����ۣ� �n^� �KL_2jZ�s���Kw҉�zz���v����Uɣ���<�v���W��=�2Z3��U�T\�l���F�5�Q-]�z	���p��[|)�wИ��-�ʸlL����b4��r�L8���<P1���v��d���fM�AL�`oX�i�̧�G��gє�^�ڭ1-]�,R�g��[-�굥�^d�y�/Y���ְ�f�b��x05��l�s���	�vq48Ҏ�L�x�{.f��}]��z�`
/\S�I�O9��aa%-z]�d.p8�0��ܗZ~D�t�@����!������Y`o֚�=�#�����6浐\)��<�&����\� ��1ox�:������b����K%k_=�I�+�L�I�[v���3N���E�+�Z�Ƨ%7�C5�/�x��@Z���"�ޕ�?�B���`f��!��b��7p�7��x"���qGnho�פ}���oFGe�r���� rXwSP��.�����|���ǈ8�ߟ�> ��-�y�m�l�H8?ʛ�V��?W�=�;��_׮s/�*$��}�L���>?+ۆ|0��6Zî�W���Bm�Ww_k�E���#�f�u���U~��3�  ~#�����b�Db_���i�� ���;��٪�s����+$z��6Pf^[Y�W��qx��f��[�G��jY��9�!�������q��|��;�m�KE��@��;/�olU�(qf�S���[|6θ�4Q�x%Og=���A��(�<T4J����rĳ�Y�춙�Jl�[�D������:ɮ[JY6�Ӄ�}�OH�KB]�QC�*n��Q�Á	G���l���6�5q��˯|sB�T�~�N�L�9G܁bB�>�]��r����zo��~,��0�C:ðt0�`�-�~q����ț�'����u��=��������w�KMڔF+�<^9�k�����Y��j �L��/�:��<�;��-Ī� nKqy���lQ�����b��c�߽����fT����f����K��� �0���C�eL!���t��_gs�ta���Lu�M����U��i��2�߆���4��G�n���L}�kd���}�LO�@;'�����Z��@����fר0>�~a���g� �S�:��}�2�(�+5�����u��]V��G2U��l��'!�.)�|���qM���^�P�n~W�ʳ0�B3tm�(~���/#O��O}���a��Y�n*�A���^�-�[:����}��٬�|C�o����rɊc�l�M�+{Jm{�梏��+��͎�)J����!�����x��6Dz��z\ʸLÐ�2���B���9Ӱ�ڗ��KO��]�W�|82��'���G.�/��`�܄���ά�N��U�=�6&�#��f�6�\�����3�T�o1E��Xyd$[�_��+��L��p���e�:�/��e��FV5�W,%�b�]�JssT�Aqp�2�ɔ��4Wd���@J}�"�ݔ ��(� �xb)q.�����W
S�Ǻ�0�/�*�ޢ�����L�O/����q�v/H!�Q��Լ��|������c�y7��,���_�XeP��Ӛ�ف^����a��6�p�n5�{|������fut�n�<��ȳJ#�-P�^�o���ʡ؇#��Ʌ5�lV��>��̾U�Nq�'�}c�H�@�m��T�@<��#�᝘�q�wc^uN�f^���q��^�{��=�].J޻��	G�2�#��F,\�t�!�n������*�4$���X���վ��{HUwA1p�d.5X��0��!� j&�K�%�����"�ֲW��v�ᎋ�ۮr�����y+8\��v6A�6�۾h�?%���T�b��xj��#���4wJb`�/g�T����)����@�;V7*	y����u��d vb軘NScgR�Ψ1	@�ȚW�łs�RN��69s�j�f��������N��ԽIQ�x|\{К�x��v~����� ��5�-Q:���e"�.#��;���}��<-y��(���R�;��p\��n3}չ�.���җ)2]���U�辥�2LA[����6J��J��o�P�i�;,/�.��PwMf�Kq��SwK~�d���f\����\e�����i�Dp'6�㛊���;�������o��p�dwh�����'���s)��`���"��xb\���{��e�{��Z�׾�G��l�]��[���u�d���}�"�Y���q����m��<\�:S�˛��u�5�yԞR��s6ɢ��"�u<As�27G�����R�[Eȵ>ޟ�qo�s¹��y��ǁGx׾�B�0��E���ͅT�D ��T��	�����(L�+U5f��=�kћwo���RĀ%��f���K�������1@���lԺ�-#��*v�{d��������0����zko�V�e�WX�6�`��G։?��G�L	 �l���/�"H����g�?u��ٶ�b5�#*m&�	p66-� r
�&1�Bu�d���߻$@\ `:��^�&d}�!�=�OL��P&����!��5<��Q�:x�²��-k�'騰�lKpl�^6L���KH��^d���m�E�p��E�C��7����ҳ�ǻ{�ù�]�	�{'z�$�!��{�.:a�N�5QG���A��A�h#z��{H�99�}���~}\���s�{���u���b�Vab���Q�p^�>J]B��}/���#���K�E��'�ڮ_�����(����U�ʳɯM�F9
Y����m���\ow�LLk�nW��.Y��?���}����H��o�!���r��]�@�0�w��C����X� �	?D�-hM�s9��#+���K�����S{�q�c��6S����0sӲ�vZ�+(^h�@�C~�}�4��F��������
�~��PH�r�m�� �	�}0�U��D��}��Y�5�|w��!V47fU��z���cw␷0
� ���2��k�N��������ʻ ����vԘ�鵿�Nf>m��hq���RB{58�
+9���9q�S��twẙ��xr���0��>��x�27hѴ��϶t��li��Υ�w[��p���}W]��˳���9|���kh�Ӫ��LOf��w��*��c<��-����ܛ��lb�d>e�^=�\N��9�S_�3�͖if{h�7n��s��^�8	���1���1ͪˣ���}��I4u�i��A��!o�/�p�H��NW��i�6�|1��WkD�%��T����Ͽ�!f/ ���+ɽ�F"����������N����z�)�ĝw��z�Ί����&d�B)/c������]�M���O�Z�P�
��H�G��r�����t)=��O�Y��Յ�RX�*m�����I�n/�������蠟��W�Fz��5���vqf�� �:ꁽ���B�v�'���'�O\&[��.�������gů���o��4� |By)����N��t1;%�8�L�2�(n}����)���h����/�b�/��v����m�ǣJ��e,����z�Ovc�#{��25�q�+O��{D�a-��1b+l=*�:u�e�2�[���.�k��)�ځ�"�<)Ԫd�Wgڋ��7�&��0�e{jhLޏE�"�7J^Q�(m�i�"@fU��t>�7R��'@���k��c�JB����	F�cO7�����F�����j��u�n�;�q :�z��^A�i֏^�����!�jL�ğ�~6�A}4=�Vͺ�gv	�����:&�>����T�ZJ?���~ֻ!��=_hz��b4���7�Ī�:5&�}�zy��&N�>X�b9�,���_�}��`�TS����iZ�7Bu񛖔��McOYI��BW��.�����0��q�q��YU��N��C|nY>�4�.�1���J�ڶ`�=�"��#��A�~�.Ը֕ci��o��O_�5����\�� ��?�.r�%
���s� Y,�������u�m촓���U�������L��O� x�Ϧ�q�O�|�u�Ru�v�h��G������[+�R�)�ۡL+ߥ��K�+�Z��C�(H�#�C�O��>ޏD�հ�B�έ�;;S��?<�=8�{.\k�%�#E�zt ���Ϸ�
�^��)�zx��:Ǉ�^y��"�WP���w�&�p�{�����}}����!�����w�	%��ۚ���:�\%R��Q�:{�@>舘���֐9�p�t+d�3�Q�s�E�������=��Sg����n�O"��%(4�4�RQ�FvD650
4M�"S۫nY��h��gJ�KW�����F6��n��7�<�Z��Ґ���'ٺO�Pv���f��Ʉ`�����y��Q~�H�?�ys��~�߁Y/���2I&^���J���~A&����i�>�& {1$DE����Y=�`��{d�jd����������o�jj�M�z����q���1w��W��9�
˩~����`�%,�5:6p�V�b!k0�|h<���߉S �5�n��j�yG����G�]X\�
�WwO�>�2tN ���_፣��)�{��vHV|r�w>�1b�%Q�m��m<�zD#d�����o�1�����s�1���`R�7g�՗/�Q��.���ɚZ��OTۢ�\�i�km�
��#iz�>o�~|�ַ�'r�Z�L�I����?�����
;Bp�S��`<��.M�IzBNc�
�~må��ʸ��r����:�b���;�;�~����[�$�=\ѐ���V2�H�$?ȗ�\O�����_�(yk�{��C������s���oΊe�!���[?=6]���*��^�U�sz%]�0��&�dj���4���G���O͇�No�v�oB񝁬Z��o�׫V������Swhkه~1�0��:8B�{?����[:t��?�?^�-O
2�Y�[^FW5!\��0�[@�C�� rH��\��9�[;)������|I__��Y���$��H�=��Xwg�[���_���.敕��K{r��� O�2����Z~ٲ���ą0R�9�]�~A��_G��P`̀U��]�Z��v)6L!�Ģ�H��:b��Q���Ȧ�<����׎��c�ܺ�f�� by�5l����8V(�{�\�Z���]�j0���0s�N�k�Cϼ�'��_�����[��<�o��L5����%�[<)K��1A ��oצυ�n`n,ڢgC�R�{l���j}Nč�~�&�o�gV�቉��(�S�Nt�	�~������!x�!�x��l��|��OP3.YfT��$>/�������Q%��: 9���� �"���mիG)v�@5�n��?�V�����Ϝė޶��p<*�l`ň�V��"�|��nj��$��Y@���|1?�[j+�]���������줗�Vnc��/)�Zw�5J6<�*���0<����L52 ����J���YT ��b�(K�����l���뻧�8a���������|/p˒�e��D��j6���8��z���;68��Q`%n���VL{8��e�ߦ0=���3NzJy��5��NCq�1P}\ux/l7s X�u�A���5�:(�ީ�^���U�����������6��-�ě���?�Ŋ���$?���<�T��H�/�fE)����<)���$��M\�L�*dy��%v��5�rs�(~�xz���įO������y���b]������*G��GX6�U�K��}���� ���과^Zh�ZK�
���i�������袺Yf����K���7�?iΑ�N��%�d�p�3y�� ��4q�[/[(\�[Uڮ����<1�	��
�	Ҳ�� �Oj^�'�п���#,v�,|)l[������c�μ+1�Mh[t[t�ARag^/J����_ce4��Pa�y�>-º���P5Q�s�f@;�7�CH�_���ss�����د�<��Fa$0���Q,+�O�;kL3�ϳN��tU������L�uzU�LZ	�^���B#4�~�}�:�!�P'����qrgL���tl5:r��ڳ}ґ_Hs��SC�� �<��]��K���FJ
�c�n�������5��I��[��)�t�Aʏ��^��w:�Ϙ;;W�ٰ�VDBX?[3CE�)Am�P> 4�рi�l�A���iP���Qj���Q��3Qf�.���t1�D.���|�ݼ[��DX��ߛۨ��0?������2�j̛���y=cM��ң^������:��tn��
��%�dEW���$��b�0ATqNW�����R��o��K�oZ=|8:��/Q�Gz�X�m��;q�93�Qa����(o%��+6k/�?p�D�q}q��0-ᤥ�]$�3�2� ��'Y�I�� ��Fp#��������-�Z<7���B�+ά��v|�M�p��xw�y䏇S���%��ǻ\>�r^��z�d���=�1Ag�t���6�k~�/b�-���1��+�y�H g�Bj�X��+JzA;}j�`�������6����ry�Is2o��Z�'��"H����- �u�x[��_��t���&���S�mM׫�EѸ�M�rp&�>�<�@0H�L�����m��>�*��]��?:S/.K��z8F�R����a@��"涇�n�>�7�Hٷ�Y�B��,W��h�]Ž����8P8b<�+mԹ�3e�qqg�x�/W��X��:��«�]����G>�aԗM���-@��)�����}���ɰ�W�zX[�Vx� ����{�8�5���a�N���?m�$�����=Y#�*&�V]$d�z�YYr�f��w�����._��3R�{�
�}cWJL��}Ym��?aQ�x�% g}:�:����G�XIw�
��3��k�bXR�9IO�F�}j�s��u���#�� �&u3�ڧ�2��W�o��a(@c@�F��g��k��ڦk�lp��4`��Ӯ�2_�f�8�"�Jbhw2o�I��� �͝VE�XH�/�&�~�@��w�#i��]�u����}s���sE� c�7���&hӢd7o_�e̕��G�{�C���0��}G
��EFStlx�H5f�5�k��qx�]�tP�j#`QPO���ICL)a9��[�N)�K���ْ��Z��^!��u�����i�#J1��P#	��*�G3�?N�Z7�7I�B^���#�2fXuM�R�T��I�B����U�=��EE��pC���m�;�G�a�T̡W����3�5����?5�Z�8��~�yK���E����m�z����\��ģ�O�Z]����G]�_��f>���!�Rj��J/9��=%�2כ����U=)��>3ۻ
� Ny�	j+�'w�o+�k�ߙ�H�l��ǅ�$kd��bS8�,<�IRL��o��-�Q �SC��\�ڵH�l$�U�X�����At���]�̌0�^.�)�?�Js#hH�]mL�2~��Ư��if�~���oH�x�}�����rnO������h£�QhM!Fɧ��F�p��8�j��A(ut��:8X�����^���V�h�����+���;�����Ȗ�1l�����#č���d�+�I���&��R�ۺM8�\���ef����ВFA��(s��
j�I���Q��M��������-�� �4a1k��A`�?�e�G
5�0� �y!x_;� !
ɟ֦�.8�ŷ�d�+�B"��� o[U��B �ҩ�%�?�pmyq��u�?���{��y6�y�
��_	#���_��E(ڶsI�~_c��M�.��k:]�K�#Kl����F��UR(r�=$�����;�s��g���eK2�g�c���tn:�k�G�?�AR���O�x�FZ�n �}�ŽT2��u�W?��0��6k-��,��qI�\�6G�������k6�������~��쓮&���5�K���0AT�N����'�\ۚ�O�w�����_��C��U���T-B������.+�l��_^}��ľv��c�#�Cv��B�{�Ϋ�J�U�=�.��v��Uc��	E�޿� ��[B2M�*�g�w����x�\s��䚊ο��V�����p9ﻺ��4��\|끳��_-*"9�u�*��`������q.xI8W���wt�z�2��W�ڰ��@��j��rt�yu�6�<$��`,	B�q�yXS����g&��NO�{���xD��
 ��Bᗸ���f-cM��d3�n�Zk��dFv���7Ux@yAL!^)�Y�H�V֐?&T����gD �?���4y1�W�s�Q��!�@rm��r1�&10�wNqn4��M~���lamp�oC�EGfҺq�Li7,72ϙ͹���o�*F�+��f�zds���٦x!��`���s��`Ӎ2����;03 %Q<�a��M�cg|Ô���7]l���V����R�2"y-
�%Z%o����� *I�q�$y��o�)�*PV�ڸ���I��͋mМkSC�s�E����&_�]�1��[� ��۶FSu��ˈl���3�"/�~�"+�[�Wӿ:[3=�a�0�Н�A�{��~� �U�1�MO�l@�]{ٞf*���ҍ
�aP��:�����|�(+~��@��]���aq֫[��5ڣŘ*��V�1U6�Z<�e�x�������I�|Vk=J��}��-`w�W��|��^{_$<.�Cx�@(KC{	s���ӋR���(�
�^v�l�p�U���[��:#&~���g����q�̶����F��צ����6�1��Ot\���</я2�)�O�(����`vz\�Cø~H�\�\��Ԇs	��}[l���	�{�:|��`M��_�!�� f}��)����I�B��I(��^��KN��Y�/��/����JϨ�����'%).���ɕJ���{35t� ��2�@Z���,@⪛���,���>4��]�.�]�l捶���临�Lټ��b����-z$ �E�yO�Yl��C<��vo��
^"�׫3���@�� �ck�^d�7�\%.�[rhe���[��}{#5I�!L|'�]���mO����3�cE�+�Rfˁ0��x�|����*FO�n�4?�i�j�P ����;���u���o
���	��s�x��)$��������@2�oZ͹��.�
�Jo���6Y�@���d$��/?huO/����9�ߜɏ�~�R�s�k  ��a`t@J��4� �&��w��g�.;� 3=�FBdȀ�m�`�d�@DA�/�����N�E�憗o��8�`� =�� ����K��`��ߦys����yd�W`�.��ܸ�7���(r�����(��=U��+��zg��\���B "����L��@O��xS& 9��`jD���?�<$��U�6X���h׶��w(�l�z=��r���+w�8�U�N*]B�%Vaz�t��1�_���;eVj��{�?����7�SgۀVU��6b�p�����B�sN�T�O�a���0�w���Д�i+{W�t���+ߦ
�d�å�AAFu�i�w�� [�)�p���Q�ѐ�`z�]fxA*�u�nf�6��'P.ӪD@���5��4g$���hèw!b�5�����` �,�����U��>s��	
G����h �4{~V�?zlSN5+KЋ<����QR"�Q��J4Ȭ�r-��w8��>��;�M>'�C�D,���z��`俖 ��"�^�vy|��M6��:��V�oa���@M�'F}�ʞ6�5���>�/�����֨�CY�T�@f�D2�@w�D�(H;���n-ɷ����m�0Ir��$}}�O������E:H
=R��ؕ�p�LI�e�n����>�\
�Ƈ������a���Ҿ�`y)(<(
`�q���S��r#�.8��JZ�e~M���K����3�!�>���_f�f��m90g��P9ѫ�D�S�dS��⸆W�@KJ�)9?;�Nj��F,e�;�	Ɖټ;��q�.\i���0Ax��a(�o����Ծ�P�z,v)���g��At���X����p^�jg/m��썪Z=�M��o�ߞ+�_�,)�d�9��8C��$#�����ܖ�(\���t~^���R��*��^rX�^~�K&Y��2gi8���[��ByY���kXW�A?/�j$�`�1�����n$$@��a{���nˑ��/�"}��U
x���������m����*��̊'È}��wn�]�s�@_�w}&C��]5��(��\�7�	ȗ擄ۖ�������6��Y�L�E��P��c,��|�����t���� i�H�/�R8�̇l*f�!43(s�$,=���T)r}����M]�d���M���>�۽�.F�/�Ǽ�q�v�Րc�<*)ϳ~�P��	)]?X��%n2�X��D�&_A���������ǘ�"��������a>���n�=��#�w�����X[������}h\��ޫ]6����/.��g�S�χ��s�p���sF��{\�1�T���ǙP�@����J��xN��|�K.��ڰ~]\N�G�����0��6�\�d�Sn���j\�T8�.j[�o��l�K�W��%�v@͋��{��ﺁMzʣy��8:�4��?:}�{v>X���/Ҁݵ���U���@~ץ�/� k�xb��C��]%���9:`j5b}+�8KKx\x$>���2iO��UDkF��叫��'�W��٬8��g}��S��hR��2����0b�س�|�|�qN�iZ����=3�:\�Fx5CM��^k�?50�z��n���il|����OM�]}���i��}��A
���	��p^�ՑVv|ޅc=����\O	�������|�3�i:�A�_y��O��DL;Mn���x��\�AXz�SOPۆ�㥶�ɶz��J��4щGb[�#\�&I���wڬ{��_K�)�to.�L��q�/��7�U����Y�,�Px�m�e)�*��5����ӿ*��k���}�҆W��֝�#t32�v���<}e#1�Zc���D5�9�_e�6�"ճ�s&v����� �@Nd��F[�WI����.�nZ��,�]�S�N���}�G��)w;5��ˉ���,��-��s�)ļ��>�����Wv��;��#%aH�(фp��KqH��D�uL�jk	\���zrzߠE��t}ð9Ϊ��Iƕ���`覥e>§��%=�`O ᳞�÷n��)�H�G�3��/ S���̺7<�����|�ҟ�p�ڳ<nʘb��ي�ں��X���=}7[4�A��H��M�V\$YGAO���3�p��=/P���lp2�|���釧g��̻�wQ��3��i��r'���4>��b�?�ıX�4,q��Uu�Yl�`y��4��	d歗x���&��^7WK�wu�#����W�g1�=)m��� N�&�����^��}�V��` �k��G�$���6K�IMjz������{6����*
3��T���[�j�i�l�V�}[��{	-�rw2˹n�0�E����p��e�M�f:l�r|je�O7�{)�խ<��CV��[j�zS�J���@..�L%�f"3�N��23@��2ԇ�����nV<=��+�Rr"�%ea��V�����aL��$�����H�al���ڍ74u_��<�y$�.��y����XU�6vyuB��@RO;-4�[����+��%y�҄m|���%��=	)��sLD� %k�F�2:=�CI�i��I�n-��{C@%�fҠ�]��`�4��I��iU��{�K㑯��僑�$p��%�:���f>�XX:5mF^�=E�r������`�"Ȍ\Cv���v?�K�!���ɞ�����nf	y�����G���w����!��x&y���(F3�ĝГ�&F�FX3���"��?ԭt>sB�����G�V�d�i�L��ԑR���C��|߿�&ٙH�e}}�K_W8�ժ;>�� #�0t]�I$�2���%AI3�J(|���#������,wQ&iǂR�X��:ܯ40@{�<��v�K��zy�ĝQkC%2b�A��:(� ������,��g��mV��M�W.(&��U��a�_"i8�U���:� P�1�\�~��j��o4���7kh�
�=�K��y���b��a�xI�"���p�YW�7+�Y�M�K��v"�Y�0dg�����D���f��H�}[Y��2iT�P���'9+���������l4`ť3���Q��X��R���o�{\�%穦������ĸa҆c�����W��p����}l��~��x�D�W���3�It�a�C� _���t�}���y,d� Uǈ5(��=�!�z宖�~r��j�2��:�l�-g��/��,b@���ߞ2���q`.W��]����#�
3����nƖ­���M3S�E���|�\�$7=���R/�,88&�}W�ET���f5�;��v��p��?84 ��d�/�L��kʷR��Ĳ�N-��c�Z�E�Z��/(��-h&��!0j���y!9�Ի�H rpl�E�`�����p"H��.� 4��6�W�;�H�S;Қ�� S{��"�⍌�����r�x}�z}L���T`D��ь|I�����[~AG<G9�I(d�4���?������L!��G�e�m�H�sh)L2Wf��g܁~�������or�Aq}	.�X~����삑y�nˊ����t����b�B�R����vD�D�r�(����~ϥ���~��� ���#-)��ͻ�|~u�zX�� .�R����_-�,�r�hv}$������6�mv�ڜ�<�|�W�na�pv^r(�XMKz���ܗ��5<�;lV�T�Ġ�O����ux9�� ��/�c��%T�?+�A��}_�ۋ�_��(��;9���.�7$�[3�Ȱv?AH���u=�E�&��g�a4���R��kM Q���S)��a&��&t�ȧ�"A�9�j4I��k�&ȣ�Lp+:���wl1� x� �\����
~M�n:���6f��U{<��W���p�p�;V�&�@�)�6:毯��\�`�6�( 8����Z��8)��B|�/��4���R�����|+_h�7�S�|^���x/�?('1'��c�������c�)��7�ELKV����.X��1<TJƍy�����6��do?�]qo��+=q�};�����@2P���ݗ���=����eb4D"J���Mxe1(�?^AL�	�9�e�H'�9��*j ��Qv�ɼ�	NX �:u��a2����S�Ҟ�]ۊ�Y��xd L�z��S����	4��Y�^�y�#:[C!�'�7�4<��:0's�s#�sӵ�ڰێe�C��S�t�G�S�����G*zY�Æ��E�������i��p�D�4�,!1����݋6U��U_ƛ�����Q<Ai�6���D�Rm�p~jF��[��%�~.��EC��	��K^�|-i�J��)���AM��~Ň����k��g����5mbvN�޷Sv�UוֹK����]M��Q1~���,���e\����߲�}��=MX3��ͨ8�m���W����vg��*��]�:;TV����G� �O0}�yd�6�z������۱6����v�1��-���(W]����Z��0n�>t��
v$��"RӀ���m&�Y��J׍�P�H�ZV�)����oVW{ړ�p���v�6���#�=K`sLi9��\N��m�!�|\�k���<ts�AO��t��?<^e���z�p��&�s��ÖۜF#�̼^�=%Ĭ��.!�u�ڮ��*���𬾁γ��A�pV�����-@U�i���n��DC<=�N�1��wqֳ-J�ⅼׄ�gJNl�E���.)�?��x�[j����^��S�<ŭ�^tN|Y�����?�2��7��h��r�=��18�7�H���W/|��쵤�﹐��V�rB�=a�f@��{\�zJ�aSi�V^�s���������Ĭ�ե0��R�%j�t�9kU��h�+L�?�(�{���:�;���]�H����RS�!_��@�hG�0����ߚ��(x{������o���`� ����/#��#�b=Η�v$��Gw�X���=-�
2���c�H��srCg��P+yK�<>��^�!	/�&�/E�^�w����8w�u@eyF��!��|nT�̢�g>�^��H�1��W�����#��7�#����3���J���j�G�6�����$�vfu|w�*3�p)#�E��t`A��p�ٱ��-GM����"�����to68R>���/+:���~�|Vi�[vp���=Tоx ��1*�l�[Ɖ����Ϥ��ۮ)�-������ŶxpNBL�[T�F��w,8�?�\C�n�ޮ̝T�ឍ�f�nm[���L��GxJ��w��<��e���+��aLoKWF]L<�����.E�1�@�VIg�}A �n'x=U�,�}���e���}��?)�Hc��$���OՏ�0�a�D�W'?�"���0EB��`�	�Q|���j�'J�!FU8e<(�ڽZ�f����,�3�����	�K^:uN�+Q��Y9X4�7#���ǜ�R�6\Z7�;4K�[��(%GQꔤ��Je���4L�i��S�er���~�ῌ�Z���Ԥ���	��ӽ��$f/�iEH�`b�Nǜ�b��t�nZ�b������L�59c�U ���Ьy���^�֜��Np5�ǯv���Y՗��GA(�2x_ɛ.�t�gk��M��&�b�c�Cې��[�"�	N���L�S;#�c��돟�B���~R}��ǡ� &�d2�+}99��9�l@�� �?z�w֮��_������QF��Պ���'�ws㭈���J�M��~�qSfޣHa`�Ȼh��d�S�\k����DI�'l�gWr�/���m�
 #j|�b�r5K�'��aC��4�����6�8��ߋŤ���J{Ƈ�eÞ�jMd�T��n���N*�-�""d��@�}�籘��q�랳s�b�U欱�ꌫ�	r�.%
n�03��W��b��0_�ou����w-G��+��~ک���=xDd�����I���x^�4�GY�J�Q"K/D8�`F𔔝Gi<y��J�;��L�P���Et�b�o�N;pfa�����o��{D��X�����wU�ѝ2���M�$��ۉo��c����a�$�l��y9y�кz�[��j�>�R;�	��Ҵ8c��[»R��C����	�������X��`���ɺ������������1�`����'����#Pw]co�rL��p����	��t�`� 5�T��F������,�|�D����E�u��;N�Z�r��+m{{�{�a'�--#�hx""���-�rQ$漧� SC��lU5Ώ��/L�%'��Z���3�b�#_����{����q�{�ˠu�F���"|�\"��˴�� }Q�%�W��&�_�<�߱x�F%���k�����49���F���)�$f3uڵ���DCD�v�S���Z��3|�hc�����Y����W��� �RUp��Q�I�\�-����I>*V����R�<����#kh���O��!�R��jL�@��t =�KaG��wk�15ө���Q*O�sW4����Pq�?�5�-�]K" ��Zkۻ2����π~��@߷GTz��Q��a�&�~�e�Ë�s�#��K���
��0'ǌ�9z���iQ>�'���Ym����%}1r �k�
��H�/���{_sV�{k����3n��M=���������SS���������C�J����t��qVUZ:vI�Uiy�m'���;��Iq���c�EG��[Nyʛ�v�<<�7�e0��p��b'���w̼_ō3�[�9>��ݽ_<5��I����m�����d���|�����K񕣔�a��!*�^/��0F����^�7h��Q_��j�z�\yj��wҌ)_�w�l8_]t�������=Ğ��e�����W�s���Aė����/U� ��y���?���Q�Mֶ��&�� M/�ɗ�_�y\�)7~�3�G���m��w��c����k	o�䡬��	2������g��[lt�ౝG��Qbv��qA��[�-C^�p�Spca��y9��W��
�+��g,�Z��.Ow�t�}6߾1��r)Q�`'r�;oB���}=2��^;2*B�sܲ�0�e��i~ L>�Y�b�T�k9W�m(���r�&Q4?�]�H~Uz���y��~�St�Aʌx�0��|���ٸ��Um
�<Px`��L�	������ �Xxt�!���mǱ�ܫa=&��g�<n�fE^w�FF��sG=�7�)�Zdo��]��9�8��{v�C�ג�O������D���n��3��s�گ���*,L/�[�#N��ޙ��<�}lv�b�����~�?��J��TZNW('zp_�vNkU�50���?�!g�.��\ʐg2���ޙ-��e����/S�Cɭmi�Q�.Nq!zj=�J@h�ˎ��·
#+���$P@�s���O����79I��	�㹝�����-�7r��x)ߓH�f?I/;H���=;��G�;Wc-��S|��C)`,�-6޾�8e}�5�]��8�����ovIʬI�F<s=a����{�.�6y�5s�l�Q��bյ�W��v�)��B��B	g�Q��F�6 �^K��P�O���3�LY�i8�KL����������5h��ޟ����<�&~2w��X�Wr�M+�tW7]D^�w�u���[}�����3:fF'����~�W��>��VQ�,�%�i ����l��s��6x�_�p�S|Q'X���_�P�M�?�[Sa�i����^:���ۇC���R�
(:Տ�?���p#�J9�b۷�����;c��b[sN�T2���U��Mc�-��j�8�Q��Ku
�:l�k�6��l)j/�؎��Y��-,RTe�!�i���w���_���2)��u��6�h8�5����]����x\�d�&��g/i��v�t��\:au��9�ԥY�����?�.ؽ���2��>+:"�ZC��+��״�  _Uv�x%�Us�j���0�!{Gw���S�ZjI>7Q�S��y�
��,����`A2��S��>� ��4�'`E�:�{��b����n��ps�������	%d_*�G�V(���N�w��*s�3�nU�!7��)��>�&�َ�L~XԞ���\���ܿ�:z��~��>�<�Uz^jQc�q�+Bn�[������=G��(�9���F�M-�+�>�]jM����r�R<.G�Of4Z\�.W�c_��H$��y�V���'���h,A�a.�NvBf:�\,�RG׶g�G�ލHi-�MÂڸ�E&��S��c�%Ps�����v��c4"Qf4}��e+w�����O+X��`��ͯ�"�-�%S��
��Թo�=��[���P/Re��Y�����xT���(z����ߍ_�K=��0��l�S�E�%�#���n�a��괸�����66�E����ص�i� #�i	��>��s��_��7���Xk�օ����o+��d�XT�ɐ�c�t-�7t撒�6c�IԘW�XiF�6yK��lA�z����hH�	�{�Ce�}E��V��c���������y����lK��e��
t����9"�R��-�J�����(�7���n��\tNg��<�H��@zh<�������Z�Dhk�m�����Ot���@ߙ�� A��9m�s����i;X^j���⤺�A�ћ��u&�K��-N���fg-�ZzNgfF<�c���]Sk�l�OsXI��3L���;�GΛ�C�͏/y�|.(�`r�'��[���>�9�Y��#6�>����-���a��β�x�i�.�˽u��w*r��v;��8	]w3��2���ꃟ}�"/M�w������1�,	����������JHB�+S\{G�� 8��
ߟ �@�ܝѱ�5��g�sG%��\��q��Sw���Q遨�ԅI_g̰��dRE>y\�\���Y�!�"K�?�ڟ��w�m��"|%����Q�zI��{􆤜�qc�Б���$��� ����O��XV��}5��D>$6^j{��OJBʛ���e����P@8�ݮ�8)�̓��Zc;<���?������
�3bZ�1B���bI� �Y�@n8}��1[�
��Ӂ��z;w��wR��u�!w��}�y��_Ŷd�����k�����Y������]�˰�<y���f�ɿ�X�̙p�Rr�'�8{�{�҂��:['�G�TWZj�~\��<�47�kS�Y�W��f0����_Z��G�;"�͒ʚ<�_Վ��p�n#TP���Rƒ��$��:`뀴�ڼR?�غߛ���-}��I4��2<��u���t�h��Tjٻ%���8�g<E)%���`�9�����P1&����k��$7���hwH)�#ْ�0알Iݞ$��4��/s������Y����}�}��f� ��	���*bg���\d��GU��T�,�����ց}�|-��κU��eIk{���Ҙ�\4�{�w"��!��^1^&nRuz��0]����&t%P45��y~jcٓ����=I2
�5�{+h���8�m�jJSR�@�2�0M70�nt�a|Ѽ7�Y�2O�S�����o��{��/�>!ED��ɉ����hE�ӓ�}!�U���QF/�
��S��B4َ�b��h��)�3]��Q�}>�⤺y����f�sk��x\�7W]���!�&/\�e_ܙ|t���lo+����G��
�o^K�irPq��p�U���{���ra�Aѻ�a�\D��S�q������n�0ɽ��=�J[��C�%�4K;���C��R�X#�G,�S�ͭ{��!�	瞝U�xu��Z����l��}q*FJA$a�GB������&,c���=e�����«Y�𐖿M�hΆ"R�O84L��c���kW��).���O.K#=���;J�nfz	*\�|�"�q�C?��u7Ev?ulpۿ�?�˶zf8�!�����T�3��³����M��c|��Q��+��i@�vC���IT�2%��U)L��J��y�Y�81\����U�u�ݨF����!+T7#�`�'��P-u�<ބ�O��B�ߝ�3ڴ��,*yn#�@v
�.#��K��0\�΃b��˷�S⓯�H��E��#�]mZ��pt������&�ݷ:���T���]Τ� �N��p���9�z�"�.�#���n�CSe뜏$Zlkd���q��A��G�|��a�����zI�y�M(8V 3�ӝ����uF��Q�ﬄ0���ڧ�ʚF��"�Ekb��p�~Ј���c�˦�Y�"Å7� �qF��*�����2��期[!�<�d��dB�_�1�J+�x3.���S�.�1$t�QwGv+���'Ȟ!ǯ����:�1ꤿR��)d�_���q�
jo���w�����z_��y<G�L���y��/J4�����8��h��"țue���6z������!M�?d�u\o�>LwJJ���K�t#!.]RKw���4()ݰt.�"H�����J�����}�?g�Ϲ�uιϹfgv�+���{��p<w��h���9Ş?���h�����wY��xS.h��;gX�zSH\p��!��3'����B�/o5�R	K�*�ts)�F�w��Y����a�rb�u펲���ߍ{o_b��e]�>��`����@i��D���j�;LZ�������H���q$����p�UP��x�Ki��U3��;=m>�k�j/��P�>��B�*jg�������!s�;�*�[�*ҹ6��̮�V�e���R�Q=oP�'��Ů��� �.4��[�q�-
d(E���m��Y�)l"<�Y"{�Ӓ��:3~���>�����*�5�{HeZ��q0�����Q�d1�͵r���;�7��Y��Ӏ�G����7�N���e9�N@��b� ���A8�����HL��ަ@���N�pY��	%.5o>/k�`mK�cYi��'���_�j�U�k���]��{�E�Y�mQ�.�3��Z��W򫢏���Y��Y��+84�ޒ&�\QA�w���P�&H���� �h$G½��C`3�sD�_�ղ�m�ih}?A�g�fF�J����7%`����[g%H�W��Hg3��ݣww�<�+D�<g��~�)�@d�IVͶ<!/?h[(���io
�n��^�o}ܰ�]L��$d��>/:.�w��/P���/��y���W�Ǚ������*�u�$qЄ9VEB��Xl���qOu��^5m���|�b�*�(�{j!w��Mՠ�a�A����!A���@�Q��f�3�=^A��h��*͟�?!�Q�k`V��{�ه[�b���kE��>}O��I��:,�)6_�U5��~�;+3\�����_�uît9��9�<)s)w���>��'�l�Z���~��U��֤K���S���U�Mqg�#[W��i�]~ݺ��^�`){��R�c��<Lȩ�7�� � ��8#g����oh�e��ê��Q�� נ��af�~Jh�"�JV�Q#���f<�r��;}Y�a�Rx�;�i��������\)-K� t����L�A8�i?!����c��o]	�aX\{��`��jz-��ؑ�D��-�)IC����%�~{e��}T�zd*�OO-��{q ���o�mŠJ--�m��9[�C+D�2J�Ԃt���=_h/t�d/��VjyA|��0B�%Iv����Dy�O�u(I���"~���g^F�rV� !r=�}�k���,�>]��C��<�;��9�YQ_���ǐ�������� �ݺ��=TO�}"����8@�)��=���݋��DI��}������MhO��k3�vri�GR|62�T���V*�`�΍s�PV$��L��	0��G8��JfiY��!�u�,sqE�o���ߋ���4rD����~��KX���\N�0M��ث� ��:�}�,ч�S��2�cm��0 I���`B0�����Y^��)6�yp�;<F3q��7iu_�Q�]��!wf��kf��h[>�Z@=�#]A�q5�FzzyYp��r	��a���������X�Qr�2:��aڑBX�n��?����'g��~f�8�N�� �`b���ɘ�J�TVU���˧�c��t���`�=�]��3)s�?�~)�œ�q��/F��{m{���o����>�O#j��z�p+��{*u������� �����?�M�FJ: ����7F��nI��� ��軏�sѱ�<�j������h�z�^u�Xb��t6I 4ţ����_��cE���'��+��~~�!J�M�Ow���@����c�v�`��^��W����-E|�\cq�{�j��w�q�ו4�����e�J�dt8�qd���� �-��5}���u
y�X��N�ټ�N��1O��U���n�}�bk���t����ϖ���pr纊��#����m�T�r&�s��:SqO	�b�-ꓱO�D�	�|�p�w'��,��`��"H�v����nV����U�Y*�I�V5A��+_�0y!]��c{�q$��b�� ,��4⥵�A�J�ȑO�j�o$n��$��L��y�=�H�4��T����}e���	�bU��M��d3T���D�:�,J���/���4��b�xUMΕ"��D�ev.GFb����do溊M'<�`�rU�TO/B��L��u�<�m�ܶ��y���4����&�_<)��6&�f�ǭUc��{�)�5�9��W��H��L�OW�dD�V`#:�(ԔZic�]c)9t)�7�ާ��D��P]*�x�
�p��u4n�K_v>����d����-aH~H�_���O�|F�m��7����ۯ4��y&Hg��ؔ����7p�d����J1���.�<�r!ˡ��=�D���W)mM�}�K!��?��}	
/"cL�آ._A���B"4��r�	6m�@bhHߥ�����-*�V�^�z��n.d���7�����|�y*���Ibz>����D݃������RV��%�0N���Q�_M�"�W��N �`�/�GH��A��j0�k�/������z!ih��\'�$N���j	m����c#ſ/$���(�t�[ՠ�RH��'�Ժ3�6ֽ��ʇ�z��}�|�$);\s������*t��{��?ӉI����Tux��whr:�ol�F��N��ֈ�wDɍ�d�x�;1ܧ�U�a���5I��9W��8���R1�8$xV=���ceu�t��N�sȴ��6� ��S\)6��x�Ҙ�z�d�Ŷ���Ny��,� ���u�{]�
ވ�QkV�� �zM���魯M�`_�v�S>�ذ�t4���BI��28�ѓ4e���s�+z��W(��E��_Ĩ���J�4#���a��1'zc�A��8��3�_�h������UF�"��>*?c���,^��t<�l�vOb0H��{K1�?��yY�_tH�r���I"Ph%�><r���k0L~��/>͚�a�Њ��b/�Y�!�AVٖ*"��(iI1A�T~d��J������X�Q
��N8W9w�J�y��O�	M(�ad*���:Ej�}��ղq�L�UtE�kw��>"K�����H������5.� �'�:���[��S%�A]�S����j$�W�J�ʛ8�'I����@q�e�'G5������|}�W��r�W+���`�����)j���ɭo�9S6��w n0)�2��<źh��,�u��?O�w�9_��mi���C0
�
˿�������^� �b��w���e�+�G炳��^��~�V%�!��^©��0�Ԭ��(t��DG*��׎M��`�q����8#H3��`j���e��h��1,�5I`�϶�6PH0��ܑ����^�f˄Z�:�]U�M3�C�^C��[�1�Y�X�����8�]�KP��<���n�8:K�=��&6X�;��
���t�ц4Uܳ/�g"L�L�45���jzOAA�!�mw&��X�p�����U.�Z	��EVZ���8���&�>3�"d�Ue���7Y��1qf�EF��C��W��H�����O)�����x�9��c��.P*��5:3ԮN�#�ZK��E���e���X�jЍ�C3됤n�(��V�|��g"������J���̨OTX-y��~`��zÜ!iيO&�r��g��>޲��ѾYz?�}ʏA6�C���u��G�ȵ�CR�k\�T�(�-XI.��>S'���v���CK�}ؗ����5���A��I.�)�u<J�6z��w�Kpz}@�X����,�����p�W[)�P���e˿Kz�8�������L)��Y����Eq<�o"_��$_��O�`�|xE?����6�,��S��i}��Ԇ�2�3[���(�Y}�WK��d�%�f�0������"�^-�X��˯G��+�!e˽"�cx���hN��O�WxcNB}�Ұy:7{�h�MS1��G��%~�|�Ӯ`���?&$��>Q�%%i��V�m����J�a�X얎�D��/k��Ҁ]���M�1�c��E.��o2�HX���&�
����[��$PrA����:���ηUާg�֐��@l|�w>��>἖e1��{ۘj��d��1�),\j��Ṟ���\���H��W�^h���o�k�S,^-�z���.6��zI`�����;�w�	�""y�q }�⥮߈�����[�� ?�T�����]���*��U �� [z~�A�g2EO�*�wG���JVi�!����Sͧ�,����Z�|���K����j�y��nh,.ZM��*�"2�O�����d���dʿ�Р�n�Rb��4+Q�Ys�×��#k�&�4�z����!�	$S#A�z쟵��)���!�	����k���D#ԱO������>��$�I�]�z�S��d�)	P�f����c`��$���|0�,�rZF�V��6����\M��Ôz��m{����/ɸf9(��F�x��:���f����<��=�B������`bn�Kn���'���8�P���Ls�Kx���J���ՙj{�𑪍�+?�,预p̝�vX�����C>Z�M��
��,.t���0O=���ü��W�|�<sl��ӫ��A�t򐲱�.b��9�(�}smb�s~�ɞ�0,����k��q�сW�

�0��O�O��м�I:����F��ݨ�̯���`����Z`�b�òr��	LJ�0;O�ãN)���Ae�`�����-9��^J��0�!�KiT�W���������[�6e*o�BV>L�	����B��TF�-f� 3�!�ۼ��Ʈ�6Q�U���Ja��b~3�#_���YPC�2:A���>�ڳsx�7)hN���*��!Pje�d�mXQu���a�1i����,�/�A���eT$}.�nᨢ��(�I�ތC���J��f�����g�1�w�& �L�w�gD�����E1��Q]2<'Ӥ�t����}�ɪ��{��+161�Р��A��c�M\Ќ��*�����4������;/�D�.��4Xkݡ ٝ۩�g�+8�B�8�8æ��X�Z@�R�R�<E���t�%a��{c�߰�9������$^8tE��#���I�7up��b�b���'��@��?�G�>��i���Cjdj� NY��n�OMT��Mx~��V]|��j����,�E�@�QH�EDz@7��
R����I�KU����8	�^˕E�*�����Ɋ�״�b����詭0�:B���)�)���W򇐐c����F��&�F����bC)�<��Ҥ����Q���-���q߄�=��C��ߕ}�Һx�n*�y+ɔFK*�y�M�.������a:���c�d;�^�\�Bc�T�Aس\��IRm��f*;ҘG���Ա������o�Xq2�5�ӚQv���i���'U���Q�L�*���M٬��- 6l?�������֋��'c��0ɳ^�Y��1F�}Xcp���赩�	��5KKxڶ��'��8���LP`Ǭ���4�u�q|�� _�I�r��:f&a�
<�s"��$�V����*($ȧ}�d�ž=��Ἵ�����|Գ�بwTQ���ˏ
W14��hp���IFGW�Y@[�!���!���l{�o���C1v��*���䳌x�G��'��ɏ���V��'��(X)b�ھ���8Cy�=*
�$�J��~����j��@�Dٝy��1k5c��~/�jQ��,L���STqC\���B��u� !���!�$���J�
��"�N	���m�vݫ��[g�ݑh%��1��Ym��¯!����~��!Ș�g��Ÿu>]h�`�E-*�:B���%���g?Y3�y�OZX��G�qB�H���il�
؞]
�/��`H!�:���#���t �|d:(��m���\M�4��'��8��oV���s�^�aNl+(��4;��E�n�\)-L�?�^]2��bZp�4�R'�r��雀]�-W�j���(_"�Q��7���X�»^�MS�*\c�mW�ņ�Ɣi8�c�..��^�y�K17H$�m`=�����w׶
A���^�L��'��ZI��D{�����^B��͇�e5A'�m���@4�.�趀��N��q2�	I�l�>�3�7Qk��K��]�a/�,���h�N)شzSHq�Z ~�%��2���1\�F���j	�n	�^@gkX�"F�'����S
6�2	,��P��d@3D��Ո���
�*$)������xr�q���J�^1�=�&�Ai��	�pk£{�3������Tl �N���:b���tg�%�:�ni�(��5j�l�	������O�	�.V�kz@�jHZ����+D�H[:oh��EIՍ1|�w"���D^��>+��T�H����yO_�u"���V�r�-�"JO�];�M�
_}�n����k�n-H����xK��M\3q�F�9Wq�?u��"U��u:���*�q	n�H}j�\Y�r��3��1o��/�E*s��6��:$��jz9�+��s��l��7��g��Z�6�K�byO����RAE@�ue�������J�1��i��'��{\��<�����Z/gVbg�K9�����]�����1�~ۭ�!�gh���F���L-�{4@D��,�u�7�6�j	M�=CKu12Ϯ[��	���|'������P�����8��	W\� ^y��=�d�óvn�;�A����(RJ�Q;{��M�J(���i�4��Q�)|��&�Z�ޕ��Eԭ�[��^)��I����#F�!
�%Sm�(�ӎ gϓޗҘ���J��=�P����JF�]bz���hr�ի���4J�ݫJ�.���b�o���bg��S�)����{�������G�+�j�'�9C�z!�,���I�c}������9�6��A�b~�J�C_f���{Q���)���[���O�e�Iy_�b��VX��'�
�L\Ge0t��]��&��|�|�J��R	�rCT,�UCކ��kE��Tn��Ԓ����]�@nذ��G0�T��1�3l*FX�d*��@/����;;�sUUuG탥�1�B��̵L.ߢ����$Sk	lU"�<妭Z��ݐO����6��x�?�~o���Z�2�����F�U.|�q��S\:(L,�'��M�D�tͷ���X�%O��~I����BSvG��d}�_Vb�G9�;,�Ǖ�ؓ�/(Y�}IN�=�i�YZ���&��q��9�U��F�L�bk�u�t�5���ڸ��9j�"��D��ˑ��n5!~4;P���r�!�b��{��w���;���&6��XX
�A�f�V6Z�JD�T�)�g5Y4��c����~t2K�������;��c�~�%������-�����ٵh��&F6�f�6ƻ�Y��M#��1��W�ӫ@���͠�^z_�=�tk��rj&0j����!��6
���av+��SL�K�^�1��۞:���6�s��l��رEr�Ϯ���1���	Ikzs������|�H�M��������u
�'2��B���T���x�uB�]Dg�=;�-�.��6�H渤	bw���Qixt�S�D�cbqet��ա�C%�@)�����U�T�D���~d�ZV��[W��\zz?T�m��&�1��9��2�>3}bU~�yQKg"�T��<���uvNg���5ϰ5�����[b��?� ޱNĞ�5��I��)�q�q'��(B��i%��I>��MKJ3Yy�2w��#�^9��Ƅ:˅~��Ŋ��ߴ܃�j�:U[��'2}П0̷��K
��%�;����#��m�\�??&]�����Ɉʔ��g�*5<���x����d&�,φ�/��QG�T��e�6`-��B�7�D��������!�c0?��W�#���9�콍
Ƕ���?��lY#��9�2
y��ҮѲE��.�)����d?xX�$�Ec�V�� �{�d�'Ǧ=����?¹q�'� �1��g��X|V�h+����	���GM��}����-���e�:�\��0��n�f�#i�k�k�T�ݾ�d��a��5�m���ƅ��� ї��݆�/������ŨX���������Ei�	�X��}|7O�Q;��/�"�ҿ?N�q�e��,SwH���{���=���;O=}��(���b��TbB�4�tg��2`�"@��{��|�����o�޿9�b���D�c����������}6�R���:�3鳡�.�c5�� l������+��f���8z�Z��ו5E6	�@��*��(H�h�F����5��1��>sWP�|2<��z�Y���|�/�n\���ڰ]��*̞=��X~��7[1���C��b��|h��%u}A�}6�J��P�9�u��`y���+�E����d_�wR���������!a=�����<�F�z�H��Ti�$#;Oú��R�]V#�F�oB®�t7ؚ?��:���B����Bo�M	�F�U�nb�Ƴ_��w	�T�����21��hbg��!*�����T�c�f�Qm�jK>��zw�l���	{x�Tw�X?�Ʌ����br���X�u�/Uwqt�'�G���B��І'�>�ẋ1/6>���4=�Ȇ�^n9/�,ng`#�B�� ����:�ح��{h��>[��=;}p�Z�ax�Nc1q����Ae�'uud��#uݮBx�C�)7|�ro�FO�-��W���ӯ���<�7�'"0���A�XЗ�B�n"��庻�����c(<���t�� �[�5�n�.��5la�J�V]ז������m;Հ��\왝<5@��VP#H�����Ha�+c�^��ɯ�#XG-
	=&u��GZz_Y?�"n&p�Y��y�ѿA�U[eN��SWؖS^�TN�tsB[mb���'�ޘtF�ܐJ�D<;�LD}D������[ۃ�_S��Q��C7r��O\Us��d19���P]I]���F�R���Q`N�����-���7 a����}9#Jb`�3�&�����1�h9��qΥH6�+�ksy�g�E��0�t�{$4O���I@�@H�����&�ƎQ[�ߙd�e��ib#����kG��}��-o����x:W�a���W7_^fYNY�_�se�@=���{y�L�P,�3)3�2�t5��81|��׆���Qg�����ՓJ�y/�+Dm�-�叞�0�ݓ���h�(�^AI�����GF��v�V��߲���j$��9{3�NG��Q������N?h�V�S�E--6]͉�'�)���A�P,������E|��i�$S�x��%-��8d�ʱ_�)5r�A����3�NU�u���: �9W���N�) ����ҸsE�����$U�n<ًT]��F�8�W�DPV�A�k�x�y	�.�U�&��eЮ�l��[�;�O�nsh����=��>tw�މm^_#�����Go�an��+]$�`j���Jb���� ��4I?�`�S�^�����?�1 �M-�ru���r{�L�uԊ/����b^N���,�&ق�7�������W�M����ܫ�����'5��`�6��_Q�v Љ�y��p|Ba3�G��gF�'?k��_�v�F�1�)� ^�/������s����<��f8'��1ّ9J�;��7���ʺ���PRc�u���]�����5�/�I�[��V� ����E���#{
��5��Gsx'l�����$Ve�����D�WD(��R�>r��4�`w���|�T��:���?H�� 
�c(`�V��d�j��wP��E^��'ɖ}��#��Z���#�l�ˀ��1;پ�J�X�S����Pq(O�YÎ�k0�IG����j�����tj��0�[�L`��D�#c/���8�ٌ�Hp���@��Tʜ�Ts? %�0�jL�]t+����P��������A3�ߵ{���)�:FD� ho9vƢ���p^��"��/�V���F�mI���gu���!��YP�l��-�qȳlU+�z�H�6�0��]���*n�bh��~�AMB��|�|	�]%��Ⱥ�p��[�X���\�)F�Be[�fB#u9A��zIK�w6��*e����^K��j0L��{L��I�=�pa=볅[6_�5�z�#A�����3��"a�7�C�o�#^��������QV�r�Qp>
O�jڄ��y��g�^ş�#��y�y�v~Ț��ly�/C��dS�J9��cb�H�p`U�zi��
�hEfm_r�A_v�V���|
�gЅ��к�N�=~j��D���Fh����py�<�^�˹mt�~D�q#FMlmÆ�Ō�4��)�t�Qp`/r�h�T�v��"Ȏ!n�����Z[#�m3Aؔ�q����+�ݼ���u�
��l�<��u��9}#�B�GiET 
�7�c+�{��L/���P���q�����Z/׭Ŧ��
�s�h��!;�>#oܒV��Ac�j�{��(K����]������6��K/ꪯ˳]��������G�$���Z�ܑ𺵵+��B�{K[�h)�H����%�{ޥ���C�� �v䚯qΟ�fW	3����a����c���_��-�/����G-�g&Ly	�#�O�j��=��g��P����&[��no��W8f�&����{�PD��x�� @L3ȉpg�������U�;�ρZL��΅P�y(��>��|:�|� �X�~�TDI}�/ng��V!t��+ϛ����n�4 �
?//<w0��ͼd�/�ha�J.n�Bd����� "�S�� ���'��P��� �!�_L���}\Ũ�Xp<�&��|�O8�[]���N�Z;jK����BO!�JUXf��ih?`�e ��_�Y�9,X�M�6~TBl�4��������yR�=�t�}�?H�A���)����n)\�0�p�_5�b�+Sm��]��l/2�d^"}�ڷ�?��q�c�u���2j��}���{�{Iц+
�/�ʃag�v#��8_�x$���𻢮���YC�/���|S�6�\�왽�qR�%.E<����4\q�u�E0�'�T�[	��Q���l�n�� �]�e��J�����.s@�${2u���E���o1���^]�Ucfq�h5��|�]o4�Pj���7�L�����7,���aq,���(��#��p@KK�~���	b�9��z��L�L�����d�qey+W�4yס�l�t�=��3�(�~���UP�t<L�TЙ�_������b�]��*����=����Q��;��016,F���SX�� ��J=;��w�Ö́�@����eoxo��ɇ3���
������M;j¨x&�]���i�S+5�%��f��H �~�*rq/�4�lK���>2�G)d��B�UTp�����>b��@O�2j�&
����%��h�}��:=�M�j���Sz�"����,��$,�m'��Օ�03�kG�]��4���S�	'}�{K��s�������y3�=&��EOQ�,d�grE�b{�6CC�k�%=��{Vuҧ�p�Sځ�cM�.^+����/� I��_���p`h���r���p��-=��8b�3� ݏi��s�����뱰��H��J�Z�ٙAMhѶ�$�1R�������2�2��/>ԃ�K]аIp"Q(GH� �7���ܴ[�جMn�.w�]�߳u�,�ն#-���^����h�~yl��GG�
�	D��h�x�a��I8��Z(�Od:���~�~��E�t�������yGD9?bD�W��.�������_Z>��_2=?�}��r>�d�J�*v���ŉЦZ��EW���J�J�)ߦb�4R0��IU�0�L2e�y�n%	勈n�{���_À�,��-]J��|pEl��t�=Z(�T'��������3�ޗ?L+|���Gp���섶Q�d�#�E5>C��8�Ƶ���A>@�)c���H�u9��Z�qe�4���̯7��oRt���k��eDH�%4g�)U�4�:K�$h5���XB7ⲹ�>Q���w�h���`�����P��.+
��B���T�/��5O2�N��
aL R�pgC2��_y������s�QU��x�Wӧ��C��~�²E�[H��`q�	�(�Ie4��_~�T�O)��X�s��<��l̦����A�P��3���L�s9}Z[t��[3�u@���vH C/�º��
$/����n �#�W��j�>���Vh<�ؓ�&����d�� ;�;M��5��:��W+|{M�^w>�� ���ʺ��bt�\~s�g����K��!u�BZ?�U��fN��喨��V9�5��Օ��{2��u:���"B�.����/����d�-<�����0��W)�쓰a��,ϸt����l��_�����q�8���u���$mA`<��y�HeAM���
�E����������D�x�K(��A���a�^fNF�J��0�b��U�Y��hC���c|8���*��=;�6��T�B���O=�;,FK�<Y���A�g��N�����[��H�uaT"_P���4�Q��Rkع&"����V�e��O�v�����~��74fN8��jĦ+�%U&����r l�����U�+[5Wa�9T��ƾ��zm�{��YK%�/��L������e?Ee�C[�O��"���^��ݤ�_V��4vv������to�Ю�Z�2m�c��Q�(�"�/s.$6G(�)�P�\�E-\Q��b�P6D���m�N�2�����u^�0)]��-{ a��~�ؐ�)�t�>>��#d�����;�6<Qbc�l���T��-�x�%���@Kǣ>k�=�޾K:��~�܋��>C�G�Y)[�$,�=Gd�T�����ǥL��7?�c}D�؀��u���2�a�ū�C�/RTh0���|�B�.P�v�,��S�Ґ���O[��	�}��n��dOkxۦ�T�Q�"H4p�5
1"o�es-���cU�)��J07��%�ShXŻ:�����7\��8��"�%�]0#m�;��m�a٥+g�DJ����.�#JL�F��"��Pw��2��R)�_�8���l�L�e�Q��C�9I+Z�A��Hdt���]��R�jZ�n�GF:���,���&�����D�{]D���,����yכ/�X�db���_4V𪚸PE��k�DEB�PNb/ApPB�v~���x���Q���P�"*z(�[wVf��j�"��y?!���$n�8.-�f7,3d�ū�Ax�,y�G���1��"#����撛�-b��/7C�}���I�B���I�iVb.����oi����r�E��A���0A��r"�ӹ:k��SNS&n@���ұ�8�-.�&="��oP�~H���hfm�қ�_	 ��9�:���;�(Z1vvMW:�g�m����E=��;`����΋�9�h��$κWUd���w,1ܶ��{ϲk�Vq86�Hq��.~�9�H�>q�`���c|�%u5X�)��'ρ'/k���$��}�]��ڽ1"	k����r}��9�.+�bӡ�q: ��YGN���2;�ۍA���(SN�+�P���z�㿅"���&_D\���R���q�>2�P4�?S��#������ �����v�g �6��jTZ]�m^�u98ZIfX/J�J��֦���u���kP��<�5��%�m�����&M�6�!�h�ц�����v�輕�jhs��Շ,y�;�Ӿ�َ�?�E�E��?����l���\�i���A�}l�����x�@2��T��W4�Qd�g�<sל޾[	\��]�o:D�XQ�m&ȫ涩(�N+l�p����A�ϱ��ڜ����E�W���\���OY���.{n����\�F������lC�Ug��Xgd����s���X,ȃ��Y_�g�9�#�/��5&,��<�6���=~=F��5V�Q�&���߱s{g�b���O�RZX���	��3~���� 3����V���/��d,����� �`-��������?��E����ר��qs2�G�+�}�������W��>ъ#�M��h5NN+�BϠA��:ʼ��A�VyJ�߆�f�?��fg7 S������3Y�? ��ǈ7�'Sd���ů��HD|+�$"�JF���]U�brR#�����s��"[Z6@�)#ǭ�7�2t���E"�=�~��)�J4��7�� ���K�qD����}<穡���W!��v"k����x1���Օ�3u����_�g���ި���B������>\��w�κ���ʮ�#޴�oi@�ײ��ͼ�Ե�1���3�K(x�c��RT�_]m74�3e����<��<	��x��t�Q�U�g˹٣3�tI��՚�u�n���t��Wʝ���!�#s}7��Fi�:R�$`1;д]?3o��"�A*t���Ms���Q��'�M�횆��ǿQnt�M��oy_���9���l�K���:�ǝ+ST4oYR���v|*P�Auf�[���fSs�iշ\Q=v�NAފ�����?.��S;�su&�3�{��I�y/;*WӮ}��7���5�"�%����}��a����Y��a�ڊ��f�A�vM�;����>h�E�������<�P�ڛY�ٕ \э��U����*D��چu'|}8Z����u��y��qj��t	VMQվ阩��v΢=&_��M���L��J�m�X�t�
F,?U�벿(1����N�aV�~V+�����^�{��'Cc����;��CE�lU�y�qk������kÙ�AH;�`-`C^b/��A޾-�ŒE��_�87���l ����Jd�wB&Hd��3�I�ti��c�^�S��nȚE����)�M4RA��<)"\�~4�S�lu�G;��������̨�J�/Φ����WV�A�jm�<9�vq�P7���(8*��wYTD���@�m�K;��ڝڮ�q�U�Ԛr{�-� u���x��6\�a�{�}����eA��>���݉�#�w'ȿ&Wwh�tXb[�5X��SzYv�I3TY���d�D��f
r�y���[~�x�|x{ ��~�t��k7��.�� �XG��i�F�y����|˕ћs3�_[`:�[��up�sf���a*/c(��?ذ!8�O��(�Cgj�-�˵f}ʆ��b�����W����&�~�n��.���n�`�S����^�e��-�j�����@Ea���Mz���A��/�/C-�u�g��!L�"�)�UG���a���BI\IR���A}�"�mJ0�5�OG+�3���d�}m���њg��צq9�Ċ�]��}Z���J����G��+�Y C��b}�H���$#̀��NA?o���#����DJ��|�Ϥ����^В���g���O	¬lU���L�i ��ɐo�e�B�/>k*�tg(	]}��*XZ�ޓ��Nߴ���m{�ɼ�����c�z���o�fʾtV{�|�*�v>G�e�T��t����=��58�&�8�WS���j�Л��*����s�7Z�;�V��t��_7�2Z�m�^���1�H�~����e<eb��ʥL�*�Y�}G�6�(�6vS�X�]2�V�1�M�W���.��g���ҿ���m/pi���1�;����&�F��I7���ԋ�$ t�M��
x!G�T�����胇K�xm�_�����͐���EP��@3�fws�&�K�<�m����tD��Ws�j�<����z�`�7�{	>��{۞�
֙�*M7�~�9�spR�T�gP>�+漊M��%�D>���3�Y�֤�>݋�r�ٿe����Ԁ�T\���ؙ�>]��z}o����gQ�e�9�«�]R��x�>G��,�hY6o����u�4i~�����3��[2�#�e&��Jn����g�Z�R�"
!�R�����G4��gE*d�	l9�������Zx�.�
i���qTh�_�o�6��z��xUMV��\�e����� ˕[�kb�mƞ4� �n�I4 ��m�2ܧ�Y��R���	�I��ƻ���M�ޜ$I��YW3�_��E��abA��'۠̇F���:��5��`��yl�����g�"�<��
-U�Ng;�MF��w����&%�)ˈ��O��_��r�0�/��v)X,�2�޾��%�	�[q�aC0ôA��;��ݡ-�S
�_����K��"u���y���@M2#+�:�B�>�O�<��GZ���j���'�Q8F3�mr�r�tZn���2���
W]+��[|S���7�Od=L��`m�w��f�,ҭ��6����WI0��<P�y�_�Þ�&C��Z�v�oW���/-�;�(N/��������F�����YF瑞T�t��� �J�[U�к�>�뇫���ē��n�γ�~�냄�	��G4�ף_cTO��/�΍��;�LG3?�vA�G�2������W�W���u(��� }�_*�s(դ�I��k����$���4�����;
�Ɖ��E�U&�X�x8�=��^Z�K��4�����>6��gE��K�V9E�Q����'c+货*���b����=�����R�(����o.�6�=�&��2��m料RȽ$c�����1�A�e�2��$w3+2�������s������}^����יc�i����Ҧ��y;��v��P|�.��rM5��s9	�Zfg��Xd��߹��2�tN�5sդ���͛��=�鈒[��K"1��[��f��>�ʻ�b�lv(��'�su��g�B�,��3>)Q�Z0�@����F�hK�px�+�͋"z�e��5�؆�8�b����&�vT�Ϣ�y�
爟 <�l�'�jm�h�q��p�:xjSa)��Ϊѓ��<?�Z�.�᠏ؽ\���3��'i�"�쪭}^����w��G�t��*�=h�T�}_�--	Z��mU��E�z���;�\"JH]0�(Smrl�5�t�����0��(�ʛj��(;U}�Bs�T�{��3!�f� ��M��'A�J	kmp��F[�hDVkM�����,&�\��ʭ�5`��k%���u�Q�::�N�R���X��a��k��%=X5�~h]�������O��DE��m:��7B �9W��%��}��B�]�`�O@]Y1���$����|_p��B�d���3�wv���� �$tt �\���s<^�1d4*�	1R����tq�[�	��6�x��OI=�b��{�`�U��Z��&�α�T�X�"�f�^2�%Y;W�Xt�������[�?�4�ʒ*�So�sn��8����k*��N��H���nbfqq�곔�~u�j��j��$�����&� ���Wօ��K�7�>���Ϡ\xy������U�����+�+Y���;#��1��S<��Ĭyױ���U���w��y:IB=l+#Y�s.ܚl��
�/�pǨ-tKNo]�*��x���:��c��^�m^)f`e�~�}5�lm`�(���?W�%Pc%5KP�}G[.*���	`��^�w"���ck���'�A��6�A����O�e�,4=�)D� k��;� ��T͞c�)6��V����� `,Y��;��ju^�a|X�Lө6��G�{ΰN�BфbalA��z��m�G�/$�0��'G\\�䃉;�����c��{����2�޹�i�d�-9\�o�RcD��g~e�{+�͗��ͼV{��}2�5U��QJ�po���˃3��� .�(���D%�U_Ņ_#]0gD���ln	��[K�k��(��U�m��]i3��-�&����{���r��8WQ��+�G�����pZt4��x<����.e�)����5�7�c��1�>�������-v,�.�NR7�B���z~�XuG�~��eI:�l�r&��Tݍ�FRϸ+�٥�� �㰕Ɩ��߹�P��什�}��y��b�Z��g�z��)ﳄK�#�D��GL�d��\�B�0��ذ, �f�FyGAr�r��ԯZ AT�r�#d�r���&�A��笚�?ʺB�u��rb��7����m�=Ř�B6��Z�r��mԺ�d�ŨIB��Ԡ%�Ff�}� !��:���H��i�P��n�_y]����*1��jQ>?SSE߮+I��y]ʀS+Vm�C
�aT��L��y-��#��H�]P���<ղ�gI�܅������qWOP{��=8���X���k�4`U����ȯ�ȧP��y�'�V��1����#�����lVi�"옿6�s=u��J����Og#GX�(m���o�s�/ =ģㇳ���ٿi*I���X�MJ:B�'%�-�e���G�k~�����zV2��k䭸7�4��;_�:�z����ğ�w|U���u}�������Vs�`�&�>�&\���F��n�k�3�x���f�(���J��^���MܶK���p��es�����`��`K��JG�bx�8�z f�+�woƬ����:�MZ���]v�o�܏�ע���D|=:V���b���.j��;�8�-�|�D	Sn��p��7��v�̖z�R�B�NF��U�|��hI�1�\�;���M\�l<9&>R�P\�e�X�yb�Un#m���4��壆
Q��*e��9��6g��X��\�S�l(�ƃ�����r����y����GBy�{X��Ͽ�0Wz�n��-Y�L�����)�?�R�	�^g�M ��縣RN�.���?Zq�g��#�Y��?��[���jnR�Щ�'!{���ȓn_z{�g8kb�}��>�2xc�bJ�����<_�E�w�����~�.R-V��bW�JtɌ��;ma�-�%WyT
���[ d��$0���xd�B��k R���.y}�}��=-4��UiW��Þ�4F=�?.���TφJ��^�?��.a�3����Vx�?rY�1�L�wuz�G Qyt �/.6�5ez�K����mq�|Q#oM�_����iL���������5Rʈr�ē������z~r��
��3f�8{p�W�+M��pYx��/��!�=F���}�9�]���9��PG=P~��0�A��c��Mp�vj�8O�:D���&��	G��5�3	��J����׈8�����i��i:���؎�Z TH�zpB��4���������^�~��8c�sA�?�h���~���ː��䍺x�e�@(��n=Jn����G�UTmi.������|��`�0b8�b�(`:4GTG�Q���W�ɋDOw����8���d�0Q�H��W��E�f]��,9��&�Y[��1/V<�<}2!9�U��u r��fv��@�i{���	Q
پf��hSv%��p����	�l�VbPeWzpF��!��T����:������CS��o��2�4&5���o7��d�9%w[~d��W*�	�pAO����y	#��t��W�O��� �ʩ�)>��~37��Eq�� z:�"̊Y^O�wڪh�_��w� ��I��B�?�)��;Y�
�$&"έ��ϩ������a��"���=��.��w�֪TP���d�������F�(D1�����'���ܕ,����&(�1��v��"7vhB+���{���U��QΩ�m��A��{/�z*�*�����ۚЀ[��ڦ�g��Ġ�����K	�m���2WE��K_c�
pf�}���Fa"G��Km}���|�{T���R�(AWn*4��1���Ka�7
��Dֶ��d�[Eq�ڈw>QX������x��0:I���~�U�C���L����"�oެWp�S0�kD�t���<��]�E����Ifb-�ұ_���o`�[�Z_s�-���\�=�q���=^���8�^
S�u|�?�v&��G9"���U����CuN=�����`A�s�Zl�r�1Z�z�7}��� �sl�Go��rGq�6����j�5�p|���<��@Ķ��,0Ϗ>s�n{eB�=|��g�>�ҹ[}��`�bO�xƔ���/{&�ܼh�B��LF�����,�r0��E6���d˩��k���� ϒ7F�f�r��֕��$�H`9~��U�Ҡ�Qҩ�{ �v��ʭx�m�3��M���FR^�OV�z�y�z�~�Fs�k�Q̕����T�GyU�j`TcY˵<pv��P��K	����훸�O���(�JԬ�dL9`,b9�5�i��%:�U�"x����u��$+a~�Ë{D܃��\ߙ���Gx�@^�B�{]o�+��e�#s�(���Kڲ��:O�\O@�ge`���؅��\��}��;�G.��_:B���"�����m�J����x���- 5?Sj-�����AB v�S�����g�o�&S�RbR5��^V �\�J֟�8��җ�;�;}Ȍ�ţp@�̪�������jclj������Je�7}�2�opn<�Й�fE���L,ޥk���|�+�r�O)��.�)��NS�W/��0�{�HV�[���5G�����G��J���5wTW�.�1Y!׸4���Hp��`PËy����տ��]`>ȝV��Ey��JtA�U�\Q
����&>���m^$��K�ӕ�Gyk%�L-O��J�Si��x�~��щ��w��ţ���k�]�{~�wٺ�5ޕ��^IE|;a�銳�OU����ױ�F���zH���Q�y��R7�Y�G��y��R���rπ���������=�K�ȷn�.mZ����u-�|[�{R��;0��?�U��+�p���֮$���o��G5Aq
(�`T�X7�,��}ws�C��w�ɭ\�l����8���hֵs���fg�&аN��E���L�.�gοП3���W0`2ȎJxx�����AN�!1�f`)�B3BE��1�-Nl�9�za>�U�]kM�
��4�@�l6'����ݠ���&��W)��a�^���l�����x�>0]�	���\[�HѮv_��-!slu�]�K��Y\	���~�P�%�d<�cy�@-�$�>R$D��]�?�И�p��{}T �P󄛾|ؙ�+�%;ˣߪ�@>k�����[�+���s������D&_&V�5��4��ր:T�Q\-#��h�L�1���׷o#_��y����}	-����ؓ��sg��ox�;����3փ�z�o��>`�e�a���-�٤m6G��=���Ut_���H�kF��ؤ�rJq7U�SM�E�Ėۯ��f�}�z�ł��{aF3n��#+K�vr���-��_L`M�ȅ�禁�~����PK   V�X+���q6 X6 /   images/d8919090-1cba-41eb-9d62-14d110867e7b.png %@ڿ�PNG

   IHDR   �     ;��   	pHYs  �  ��+  ��IDATx�ܽg��y%�V�0ӓ#�03�9G"�@0��H��$˔-��k{���w���?���l�eK�%J�$R�A 	"gr��{R箪{�[�@K���������;�y���O�7�l���a����7?�_��sw��{>�@<�խ�ہ ��p6���+l�^�&�����Ŀc9���/�X"�˛v$5��d��P��O%_�8��y�\ʓg<#��Ǘ�y\���g�~_��f��?q���f�o����x-���i���6_�����g�i#���P޾���l ڛ�9�I���o�+�����y���&M�e�*sV�/�?k'}����<>��~�2J=V$��c��_�t���X?~m����}�_��?��W�\>�Ϛ��۝���v>?n�y+kZ��Ӱ�i��l>m
~Xy���vд�e��6,ôMò�1���sY/�aZf7�,�lar1ø��o��/!�#^3k���@�>�-����%`�,�^��/b�^nq�^���}kv~���x�=��\��0�o����z'��4����kp�נ]0z-^��	1�v�m�6���MKl�����m�e������ß�8�ao���o�~x0n��all_�W���[��h��c<�搊�ҁ��
`4���8K�L�_fZ��	Y+�%��c0�/"A_q6`f^�֏_�Ɵ��S����Z���{B�����5K$$�Ɉ����[sYSr����_0�6L��_5��P�brJ8B�Ia��#��/"RgP=zg
q�t&�cL���q��~�8�q��Ka��$q���@{'���:��u�x�x����}��������^W�s�c��/���<����^���o�Ɲ6ۊ,�����+���z���{��v �oS���C�>����m���xG���w��A��'� ��ȋǏ~yL�y�@�	���c��$��X�;����q�`�z. ���'�U�|4d���k�~����X0
茟Kt��;k� &��g�<:��ὸ�N��1�},�ݲ�: *n��w 29,�L�˟|׷I r�k�Kl�~P�7���]�����31����	sǲvϳA&�6�kM�!��/�����9���s��`K�
�w�H'���u�|������3���x|���(��t���[ ��q�P[�5ms.�氎W[�8���lF�ě��o\珠�̽�����>	?� k���C7��O��P�xN�1�����4��np��׉�Il,:i�D^�^�	��Ce�(a��������̉3���@0�+˴]��r���e����Jvo��g؆c[���G����L���j-p��p�-�!�A�
�9&
����sMG�Y.�3��/����+S�uq��g�.0
�2��\`y��Y��ĵ�e��;ƞ��Sq�B����2i}]q ��9,�L>��Þ1���d�4�bJ(���1	��3קF�~��ί���~�ޡ�X��ӹ�b|��$֒��*[�an,+���5������|�>e�a����!s�u�郱j>��^0k(]��,~s`2�L�La�<�fXg�r_�
L � �l��Vv�+��O�f�L��6��`�˝�뤃�!�W�^�FM-�a8�(0(X�����������{�), ��m"�B��g�
Sh��_�P,�U!���23���������g>�+��1��^�̀�rxsI|�rP1v m|"�l;^*R���o�w���0�9P@ҙ����<����֋�,3@e%�I��s�X���Hڇ+���@��1�d
�px�cLL�#l݉3���s� �2 �`�3�wM�#��� �0Q�/?X� *�d9�0M��N{T��Ú�p�m��l�WY�n�!��qAm�� �ۼ�J5�c���'Gr�>��e(}����Yd\�j⬻4&������L��t�B�����~�a�r�,�-�q��<�2���X'Z(S�^�W���],|�E%��D`I�7=Y�be��E?�����lO��~�3�R?n���}M�&=�/��Ob�(DGVPg&�F��X��@
)�<6���<�:=�C��p28����*|++�y�0�l���7l�����/Ra̿{
�c�,���L��N��añ��-�����G���s�wm����2�	����cb�*��^�=2���*��r l��FAp\���X�Z|X����..���xd�4�R�8���D��%D��$�6e,�y��l��1��,㜙:y�M@=Ͻ+uX�h���l�o�y�@  ��tÛ)5<�z.`��4@��8��LB�iNhMy����H�HB�bP�Oz{{��@�����#���~o��8ޗ��T�I�\?�סy��թ�e��S r��w��x'D�C��A�G��
㻽2��^��ݯ�iuȣ�{��I�x� C��<.-�0�d(ל�Xw4��o������Ͱ���_u$
H���8Pl����8GN�|X�E�����o4�'�U�h�|��8E��hT��-�DJ�����r��%���/%���O�pp�p1��U� G�dC�V1��1M:�"�^z��.��L����O�^�0p�RɄ��J�~�S��a�òl�"4x�Lkl�*4>4)�����n9|�>vVn�uHI�$	G�e41j��:̢���$ԃt�p�Ga���T���c��P�X��i��Jo�n�m�&���Ý�� ����;BڍI����S�8w�P&<>")����A
ޘm��OjWA�y~����s�>��@�	�$�BK3
�E�M��u+��ˬ�i9�M�!�Xâ�f��5ˤ����<wQv��H���?j)��W�'�>p��i��׺7 [ V�9�JauNQ�g��%h��<�j�s+)���N�=>"���g�|L.�+��5226&cc#��������bQ�<��9v�|�_^��/K<9*�X4X@'�"؂fӀe��� ��ftյC�萉x�eO�t�x�n��+�vV�N�ug����,
�� ��|Ѽk������G���=a;_pP�ym���a��Zjw�ǹ�D@w=�R!k�S����h�3���ӓ��<��'�G�B��dhpP::aa�RRR"�ٴ�j��/E�e�fQ��Z�$����r�s@z�ú�3p��T�ɓ���G����qT�ՠ�^Ú����1�����\�l�<��2��I�����
�HQ��T*!�!�\���:Y�|�4Mk�����~����cyX�bu�rt��ry�k2�
�� [&\s��\3aV\3h��O����iw�s"Xy����a]w ｗ!�] �]^�]�|b[�,$�Ft>����Ї �����~�,	˗��)Ol�ո\�ňF��5� �:�J 
��2$1,�4��Jyt�RT�7�= ���$ϟ�����q�4�p���"��)m�kɩ��E} MR��Q�%��x�y��g���T��:%>0��r >��� �<yh&��IՒ��x��	ih�-�������%��I
,@���J�n����ʻ�8����tuK���,g�3�rw�~bB �S��Lù��~�w�nS���}�]Q'�j����x��ѯމ?�jA'Bܤ����d@M �m�Y0�o��1��t���R�>����Ѓ�����II������`<S��r���X���%`�ἍI��ɲd0<��ޡq�|3΀��Q�ɧ�{������ը9^�[�0����-R�TD��2��ACc�mttt���Y��f!��+���O6�[bl\=���))���6�ŋ���1�%	9.�Gׄz��8�E]k���"=n|���TUMx���a�����ٮ�n;����uK�g�s��*L��s���bH�t�6q��@ES,Ƅ�r��7�b�{���;�߲��pq�C3��\s��@�g���;�����v ȆS��~h\S�W�vt2M�9�L^�ǎ��R?u��_��Z�󐌍d@��c�-����Hag�lv��PçJ�'tYq)*��2c�f�Y�h��t��i ��p_�~��y��z�n��觐Ws�322���e����h�L9s��JQY���>\���.�bl�r�\���R!�li�ˍ�[n���L��d�B��`RL��u�?���Kw�։�;��r���Gv2��V�t��"�pڮZ�Yໜ���<&�eL}͞0;Ca0�,#>��r���M��JmeXn]����@GFF4��������h�<~� P���SK�Hb|P�++d��yr��5�W�D��N����	`��y]ٖ�&V�:��b? /5�e��<�aRrh������ ��9%� `�����ޠziIRm�V��?�%--�pa�T�J�C���bx�q3q�N��3����:u�0���x�0�8Ὃ|���q������g"
`��,h7$��4<�6��۪x���>������+$�E��]�����Y��=�b�� ��࿃tzrt�M)
zd���26��II�e||\���!"��I�L�9���jC�)`J��Q8i�2�hQ�4L�����r��[���a\C_O���X�rԐH�>�t"�~�_�`�PqHB>KfL�*��K_<��zn�A&��)��O���(�������1M�?q�Kk"�kgevK#�Z,}�qtdDJ�K�2��p�<N�	 {���u���lMk@� ��hJI���g����>���l&syGK2HI�Ĳ[���y�  V�N���aH���&�\�u�1��k5.G������^�S͐�[jڹ�l7 �Xs}l�D~���1��?�+؝$��;,ٔ%��c�S���0�V�cQJZ����B�%��F{�'wi1%g��g( ��^��W���|)\G�Ú#f]�'g[�#@n��37��4�L$c��46��%��y,���h��!x�����(�x�?��<4c.d�(&�<V���w���|V&�u��6��^𶕟ȩ�x/Nt,����7rM�臷�q���]ƪ��^MS�F3�Ҵ��=0����d����LjE�_'�r���\5��A����(͞ǫ�U��M�G� ��\�C��"�'��CeKM�ݓnrbf^W[:9U��
�Y5�x�7`h4�k|L����}z���@(�Xl��0ːf��9f�e{�5�^��f��B0���1�D�`>KS{�3����,{��9L\�1,�յ*�ѠhYT������TB�l�kD��9z[9]A���$�����c�[@ɄD5N�eJ(�o?z�qJ`
�C�Ƅ<n���j0�|'�U�L�Oi��,�g�B��"��T�'�Nb�3j�`�`�Q/�׏�Dc�RQV7����9NR��!u}F0I"�PD��1a]}}�70$�|J�K�2ɐI��%gsXpL�c,Bѐ$���@�cJI��:-� �_H��Zs"��QMib�X4�(�ǆ�!�-��Ӵ�i-;b�2s:NSk��aD�C��(�{�S-�����7	'��;y`��1o
��ܶ��ț�LF#��|�҉26�+-�Ϻ��	9�V�}0^mx^����|��3����f�懥-7mS(+�N�b6޴�����d�Qt΂Xu꣌,A���[�b�0iQ)LCEm���TȔI�RUQ	/) %�Q	��������:�_�Hč~{5?f�mwD'+���gs����Bc�S5�RRZ��x�� ���&���[z���`L"�R�W�o_�E��;�z�N�����yY7��,pq4��o`P�ɴ����<L[@�,]�Q3��4���h8ð�S�m���� )c,�C���%:p����p�}��{����<��M�xԃ�̤s��b��h�	�~'�a��a�M�[Ӝ��;	D&�S�NT<>"�� �ϧ�@K=lө�q,��D75'��+�AQx�o�ᠮ�DjTL�b�c*�&�E�jz�̘6Y&�U˴)uRp}^e�p0���&,RV�M͢�ӈ��(l,* ��*��3�K����J�2��$ ��GF�Z��'��c�r~���ё�1���;���.M��S`~����'��L�BR� e��C�ϰ�m�a� ��!���8���`��5eN���!�L���Qs4��u/�Z�OE�ᄞ��iik���YR	i���i�>�Xt��p0�,�uB]�����q�kNCd�~�Qyq����>��Ib��O!L�u��`�p�HM�͛7���&�R��x]>}��\��,��n�Q^�jZ��j��Wى�8��q���5����u�R
А�6JIq�����ҙ����.xA���xb����S��
�� D0'����⽪*+erm��~��Ur!��=����"��14����b��y`�Or��u9�zU��u��I���3�W/�-�qL�3�Z�H��qt*cY}�mr�\�47n�'�S1��@��`�,��H%�n=��{fTO�%6A��/g�ʹ�W1N�D����r��k[��Xp�����vKFl�r��{$*�|庌���A&b7�W����&� `������2L5���LBm~yeVT�;y�cD**�ieC6G���֝T�9����A'�l�R����gU�H�Ȣy�4k_�:
�V�׋���p�
�aLp�śr��-��6��� <��x<��R3g;�/��p�Ƣa��-j̩�Bx�:̽���Jcc�L�6MJ+�e���2uR�Sׂ/2���6�j��Ue�U���L6.{L�ɼ|t�||�������owH�pKg��Z�N�.�$8%�h�u����,[�@*�b0cYSe<2���X���-]�7�T���@�1x�I�����H�X&ů&�9��X��c
��o�QVt�-'������:{�ƭvY4�Y�X��LE��Rm*e��g��'5�ϙ�Oɔ��t�[�]���!v1��j�,�~����N]<[��ҍ��6�xr,jH3�i��2��I*K����Lb0�t���{b4.ׯ^���,=��
��>�[4�"��P�V����+*Vv�e�Z�G-��͊KqY�e;)�vx<��^��֕���8~�X��-
�l�1]�_$3�̖ںz)[0_�Κ�,���.�/\���OKՔٺv�<�i�\�v[�8'>�V�O�OyR�e���s}���*+E��r9t���=��|�OACl�V�r�XrLr�rnE�O���%�!3�x����sf֐��
����)�d������;:ɴc:��r��֧1!�p_:�S/%�՚�IjP4��)��P��B2�LB�$%ZR*U��r�V����ץ��OJ*&�"�(
b<Li(�b����(�`&Ä8͍k�{��Y�|�4Ϙ&%`�*�H��
�"����]r���h�)IL��{0�4cU�%2�)ͷ,��łp�a��	�	^�X��ьSC���egS����OB0/A��ڒ��Q�s!1�F3x��9y������T��dM2k�<�9{�̞=[�7Ɍ��%Mt��y�}���/S��d�W��>�U�;����t�h��x�F�l��ةtխ8h2#�J0gE=ֈ��ƻR\\,�yb�����l�5s	X�gչb�o�q��Ln`�Q~��#y�/��_�Z�������$��S��$D�m����P��4�4� 7R䭴���a���x��ǥ�!&��^���Oj�
�8��]��.�^��.����r��	�/&�5����!g�Tq$�Y2��OC�ĢY�|�<�y�4N���1��83�;��gOa�J��s��F*)�JUqz�L���H�Dz#�3<0�Y�\�K3��O���ʔ,�f����T�z�Ձ���f�ʀ9��2��Z�Xq��0��e �*I�����r��qe
y��-�p�|i�͵q�䰀o��n�ɑݭR;�Q���&y�彃G�㓭�d�5��gi�a���$U�v�K]e�4�^ 7Z�ȷ_������'�iS��:u�\i��N-E ���,1�Ҥ��֛o�~���1�E(#R�^-�Q�
6����s`yX�@dA��s��T�����S���[������%sen�4��0Dn�0�K�w?�a)�����!&/�O�k9|⬄��RZ^#��I�d^��
&��8!�#}�/!ٺq�l\�RZ���Ȕ�Z����>yR^��~9r������S�V7I�����/tG��]����l#�;�mV@`�r���Y0=O�z��3ؗ��F��,�&Å�R�����w:&�t��_Ĭ��a,�(�s�a���4�C������FV,[*7��9�gd�`������ȡ�ޔ�I�ԖU�i�r9yᒼ��{r1�'�<� p�0M�>-�CR���m;=,��;?�3'O��yR�Cw�b]8ccc�Ҳ�8�pR>>zN^}�-ٻw�t��I�|
�T��<�<8Ņd�@ؑ+��7�Aﶊ9�+3�r0sn͸�yxY�d�����/@��d-�dŲER[?E���hH���.Vu{{�||x����^���#42\��M@���0�ĕ�xo�W*b!ٰy�,[8[�.�#���9���}�˫�yYn^���&��p�,���XJRR�XP��n� V�S� 2����i��������42��+E=N@�v�/SZ^��DO?^wL�߫�@�/�������,?�Ɵe��e|@c�51.{w����sf���ҥK�f{3�{{�?y^���+im]�@V�o�_��B��\���͠��b���w&?,� ����g���L����5��8�V�`�n��k7nʅ��vX`�f�%�4��gaeAo�J��b�O�@0�7e����fO����*`9��sB��
h�~���y9�zN�~o��F��s�5�z�u�\���=L��JxE�2bLĐD"�Ca��9��!+ΐ��Zd��F��.��*5�p�����+���k�$6��N*J�4����@�i���F��Q��(c�7B.*�ջ"a�[Zf�ޙ4i���AQ��V�������
���18�����ޞns���G�%���0k}ii��TVA5����V�`|&f�'ʄgO���dM-Ͳb�jY�v�L�ڀ��r��m9{����,Z�X��?�)���ۻ?��g�a�d$a�%��n���3�@q<����Sr��%9�z�/-1H	���$���P0�9��&�B�A"@_[�`'�a��M�hT>5�l���XpU����l 5�L�&c-إs,$銠@���w�_� v/���{T�3��<��}��>X�a���ȝL��^f̐���Ʃ�d������e2�*/�C P���[�����ƕk�M�Ҁ�r[&a$>)�U���S0F6��~%a~H�)��r��3g�ܹse������u��z��8�M�����4����qj�㨼�\*j=2{�2'���3�'�4>��ڶ[7�����5�0��a��e��`H4��F�@gй��C.]�����߱�1il� VKm����/| 7�^�%k������P����r�Z��)Ї���
�\�#����j����C�����cOä� hU�s��{�%�Sq��"�e(­�2����?�cym�Guh��sgw
W'i�	Z����O�ǌ�EJ�"`���3��՞���)�F����y�f��Jt����a@!rCY�b�<�c�4O�&L�+���K���K�ͫ��Jej�$o0��,�r��.1=#:ɱ��$��bp��<���Ol\|u�/����!�:$��8�+���E�� ��Q0��j&��h\t5Yqԉk�N�*S��X�������ȫW�Jww�� ��A@�M�$�X��QI� �]mm���{��y��g���-��:��='�/�?zO�L�.-_(�[��O_yWv�?*)�2#V*#ɬ[����76��Gb�1B����kԕ�~Q	�� '�D�{����Fwʕ@>*�3��W�|�)��^'+�=~���N�Q�p�H�V&�q-Ɲ8Ь���H�k"r��>���Q͓J�� ����`���D}0e���ò�B����0����!)���IS�z5q�d �d��`$�����e�0����seŚ��l�J)��ae�h2!c L���:qKxh�� 5y ��.�!�L\���ѷ ��!$ �k��1}#��y<gL:֝J�0KW��(��4w�L�5�q �����k�/ޏ&5>:��Ή�ue`�����zz�@ʃo���y�-r��)9z�0�F�,\�Q��'dL�O_~">E��	h`{,�9�d��5�����F��A�!,���U�R	E�:���K��RkĞ�TB�{�Ȼee�P@ѥ���e~�% B�2��Z�R��e�4�jFw��L�d�J�x1��ye颹�c�f��1�¤��<�/ˮ7�R 754B��ha�ϫ,�B�0Q��� L���n�4��<��!�p�GaZ�:��u/ldUa`TW�OTt�������4xf���J#�ЀZu�5��k��v:'�u�b5�5���z��UUV;���Y���V,�������w8k�ri�=z-�ʸzE��2�,��ݚOe|������=�x������2c�)����w��Y�l�<�u�4O���m9p�ֹ�Q�mI�	=�@ ��`9r@4
S��L+ٓ�lHޓ�2�|.��ae�V>a�#mf�o
\ZVm�;��0ә%��[>�
�9��-��o��h��iV?��L� <ff����fʣ;6Ird@:�^�J��[e��Oꪪ@�ͺ,�JO�b�%���d��������U�+�V�mx5�����%
� ���o���K�J�u0Y{{;�S���Ւը5��G�����QS�	cuS�ϛ7G�g͔��3�C-))�
 �_4��dJ�MR�q<	��/��bp@�M�"�0��5U2�c��^��E�T"�}�{��.݄��F��x�7 �My��_��Z�H�(�g�I?��`�*�����4�v@~��[�"��%Je�2������N���H�ȋ��X9�nF���,V���ӼB���d�ޓ�ts�m߳��9M�9d��"����Gw-���)o諊Ryh�:Y�r	��2V���1��pMN'O��a�nŦ��D�i����TBݔɲy����m*�����G:4�e�������DvtuˡC��Ƶ�:q��,<��z����2S�&�)���NuwvS���Sg���Bh�"������?���<8
4�E�] �n��F��#�.\и٤�u���T�544��@\ٳ��O�OQ���)?������#�>�E��p�z�W 菜8.���2w���S��b�宣w\��%����}��PL��F^�[����;��x&N�)�t6r،����0拾i�>T�����*=�Pj�.��<�25@�3 Ąg5�+�eQy���K%���ӧ$12$]�7���l@P0uTЃ�,F��`�1��*��-��m�<���ڕ�j^� (����VY�����W�>�9�����ˣ����eʔ)�.�{ ��L�U�g�y�$Z7�2a���$VR� )-)W�2<8��μ"��nܸ��mj%���<xP��٣!����Qf͚%S!�S8n)|WT���7�����
�F���{�;wN��LnS�����������c�ත u���>rDΞ:����EгQy�_����b���A�B�pKwC{�F˭��h�����lg'��/���p�}�'[8,�川���-�7
�� +l3w�M��- �Z>��T����A�q����4Y>���� &�<�R
�	����*-é��fHzb>VtB��J ������O>)5��ȭ��:�x�Mm UI�}GVy��W��7ߔ��[���[�N���� ˗/W�H��>�Db\��S߰*�c^����¤��\�azG��8��Q.�!|���fa�AM2���M��P\�F�8p@~�W���7�ʕ+(NLl ���9���.�[YE�ԡ]��XW�\���d�}/�^�|��w�zGj��d΢yR[U)۶m�#����ba�ɪ�k$�ͯȏ~��n�a��Gʐ��@�&�-g����҃��R8��p���N}�է�t|Ή��ݛ>'�m`4���-�04f�^����N*��\
t�2U���s��7��A"���T1	�ך-np�4���y&�G�eJ�4ٺ�QY�t��%���wwɵ�u�9��0�4W�oޔ�����>��i�&y���e��E:����99{��$�O��hP�144��optP=..��0���e�g!-������FX@�kfW�de�<gH§�ϣYc{yMڵk������6oެg_�`2S�v�3e�Y���˗ɔ���^70^�̓�И������w�I6n�"�@��d�@NFn\>/�ф����T�����/�DN]hӴT��k��U8=��h�Q@�6��S���=��ҍ&�my�=.�w��/۲&���Xa˝�&��;�$�g�ɩ�vv�d%���e�̩��3��h���`��Ɔ%�h����X/5<0�l�`^����R��-�7����$w�|�E9v����5j�=����o˫����jɲ����������"[\�z}���p��L��̩j������ؔE���bQ��PQK�c�ڥ|&���F�z��Ì��U
��#rNH��V9�%�J�?�Sp�s����o�*����]�^�,\�^'��AI��6�$��
)��~�C�Q��E�v K����^u����6��N6��)p\�\�)�{_�>�I��G��,��\�эE�ˤ��ޫ�n�p,����3���tcy,ӆ�3�|��Ŀ��QX�	*��\N]������@�",�����Y�S�3�o��p�����X�u5���%�	c�S|�O#���%Zv��'��kW�[�jP� (� �����:��M-�}�k���/�6L"��W_�C5y���X{����V���:��2E���'S�e�<V4�hњ���:逓P���A �5VW\ ���G���^c| .Y�W�ȟ�Ęn$�@�'%vj����U�84���?�&�ر��v{���R]U�&���n�F@����b�^܄>���c��ڗ|�1������Z|����Нu��m���[r��	��R��_V^z�]�u�X�&`�8��9��r6]xL�0���2"�d������}���z�p8�Ӕ�{c.�g�+
���O�0���H��|�$7~�W�̰,�;C>��C��]���:jjm�X��`E�@ƴ�.�Y�+�*�LX�b��m�<~���j��_�Pc?G����gX��e(����H��&лb�7Ex1�(�s"��ėCx�%�r+����\����>x�f�j�TF&O���H���8�_J�M�!�ML4�1��5��x:���(}^ϙ"[���~j�}>5�=M"M�֒�����c�o��o�T5j"�Y����LֽO�~R-�IRR^&~P>:pZ�T%Agg����}���
z�!8@����X�?��;��o���C��;����*�F0���|�e�\p��*������p�F6��?c�4u�����I*���!螬{��s�LJ����b�)Xj�`P�m�Ƕm��������R�N35��J��Z��n���x"��.�d��� �M3�ҵ��{�0�����Bh�1����N.�����~�O�q�4I�~ǰj	$l!��~p2���O&�Y�ζs��\r&���J'�b��3��+��!��x=�q�}� 	,����z�],�9uXNZ�r�6e�$h�.M��1Y{��3\A`�!houu�>� ���,ӐE���[oɲe˔�y�+M.��� x���̙�9�U� `k�̩Ӛk���"��ʱ#G5 ������x���g%�d޲���<�1�ˮ}� ����r��t�����B��'+:gpj~5�
��^!y�pЙ��M�N����q �Z�H�1��X���y�h�Iƻ��%��a)��(� ���Q���2`��lK�qh*�x�)�,��>�����T/S&O�}{ߗ���F��o~S�_�)z�<��O�vhj"XyV�ÄRw��������~h��.�/�dB������GG���d�2)��"�a8�9ܻ����	X���֡AФ���R���{e����N�j���s8�R	|j��{�T�Aǀ���P�Ift�r�Yq���r��)yj�NGˁ	*a����-�%����&�EN=�,��;�7��n�csM��Ro\�:)�)"���Z� ��&��+2�+c��#1Ǣ�݃���ι���OT}J�=������q�>Xǳ�=v=���F�d���*$�Ӭ�:yf'��h��y�u�H[��`�2s�ԤqQ�(�l�9*.
�'RU_�/%�p�h��ܤ����ݻ!v������$1:��jj�X��#��k�{���=I=1��o�&_��W��o�o���� ��s��{�B�w�F�y�M.b�g͙-7< ���۷����왳���S"�<��,�>�k~�<j�z�\�pN�S�M��
�P�����,�2rJrh�	4V:p\.�bNk���h�f�k�56w�<Y�b�����@�6���8V*�3�����xV o�g/��L�1C���/�<`0��=�\l#��KK��2��/�z�e��7%xFڙ�@���S�a��F���X~0�B���)�v�[�u��s����舮���"IvHȓ��>�]r���|�W�m����&���[�X%�U6TW6���E�+,&��{%Z��˗*���?�(��Ȭ�-�o|S����W�`&�U��Qn�.����~�&�AcJ���d�i�̙2�z��)��� �)�G����9L�]�4���m�o�٧��C�����i'�FSC�8 '�Z$7o^;t�㛧�j��]zݢ�Kd���'�X��pH�5w�h\D�IM9ޫF�SxN�5��g�n�t�<��h�_�8L.߼~K����Y'��K�[���J��ʵ �y9t�yt�cZ�r��8��KEi��Y���Q��O_�s+�0y�p�{uǵ�0�n�#���چ�)�~���-P\�'�B`��'#��q��ϧ����7/���/����{wi�}II�ݯB�b��q*�*A�rGK1D4C���P+z@e�f:��aa׮]Z��g��;v�d����@��4�I����z�Çɶm�(�;A5M��ŋ��\�xA:��d����.z`dA��$LoW�m��fih���CnƝ9k����Hgw�:K!���:��:�X�H��?�s��g��y��i'̚�"�=�ƛ��a)�XD��/���Au6��k58Kf�3^164��"Мj��&��INoh�tҷ��my�?�2"� �q��\%�%���3��c`�bY4o�V��z��,��ŋ�HQY9L;��Ј���<�������V�m��O~-9���Ĝ�tݗ�����<�ܫ;�?���k���"��N�xE�q�D�ua�p����w�����4�Vv]p�[�Jl��Ih 4M-�qvVsC�K����������Oz�B�E�h���r��Qپm�<��C
�����ghhP�C��;wV���lܰN��͒%K`c��.�k�Z��?�U����QX�4�|�<yR�6��=��}G��Q��߀�IB�'�p���D���<'���G�M"�fƌFeI�?nx%�VVTc�o����|�ݏX�AW����R�{F�<��%=,��"(0�v/����/H�:��Dc��ɝU%`ݹ��F��WV�$y�?HKe΂%��0CwDs�Ξ8"�0F/<�CN`a����RZ�"� �g�2ܝ���3�|�Y����ex��mi��=�����n� '1)�=�Gd(éY<g:<��r��n9��~i�4Ej�q�g��zθ~	Ot��s���X�W)���q����i�l��g�\�rU����d����	�Cs�X���F������s�x�y����_�9����ի��`�嚵�tcjoo���CFGG�j�l.z��p���;^L����i7�W���@xr�Sr��-ux�Ȍ�&e*2* @�'�"���K�9{�L�4U._��)�M-�b�*9�}�(�[��<�Q(����;&��N�D��LJ�2�������J��o�o�����J�uau��� �nܸIn���SWUV�B˙���\�5|2f�����ɡ��e7�P�`�-��E�)׺��g�<a�q9�.�x�30֧��|"gx��L̳���F����Ev4��H��c��i���wJ��˲�פ�_����Z����0�O����SX�Sc2i�4���ń�́��0�̉{쉧d˖-��)p��w��V �Nk��c�Ɍ��r��Yi����D����$���/X8O�F���羨ڌ�������������x��L�a(��{�ͮ��'�B�p��j����,� 0����ʪ��v�`�iZ��Gv<!M-3��kr��E5���^�d^C4L1���-�=�3�n̳F�`�����߿�����_0��Mo�G,�����+�]��Mҡa,������Bbhk��q¥�(�۷[�����������rk�M�j�l�L��sL����BO����x�d޴<���0�$��p��q���I��������e12��I�?&�K<!�Ei� 1H�^V�B���jAx�#,y�M�{�SI���>�l_x�9��E�@�X`,�P��ӧO����er]���;/�7m�}�gr��G��C[�u��S�<��#:�<���f�����:�Q+t"��і�Z�2<2� ��'��zF�f`��(X6�vMmh��=L�wt��-��E��g�\� +u�ǇNH}����ޞ��z��.+W���Vˁ�wˇ~�y�Z\SQ^���'NSFk� oO_�{~�W����?���t�?��|��_�~�lr�p,��1F�������o���m�t�"���q뺎��G�b�-3푥0�5e��s�v)��?{N~��	I%Rn�K+i8�Fy�8Ҷ>X��~�S&��r�Xj�h[i� ~�κUKe��{o�,}�-�Ӡ���r6�[����5���l�h:��� '�4 �U�SQLS�r�f39HN2�:m2�w;��EM�ѣG����?�U��}|�j��M0k=rZ���_��N,+'֭ݠ�cY��KW���ը)y���r�f����'�}��K�c�C7�4ˍ������;'y8��Ʃ�jҘ������� K���!@�>�]�c������A�oٴ�|H��b� ���2wYVA3��ʁ�x����w��]��?�se-�z�X����� ���7����jJ��p��G}$���JS�\������fA���gd}]�<��Cr�J������˩�@��ѭe!��O9m��ɏLӼ����Fڳ��)4-�%!y���r��Y�:�Z]�^.���w6^X�@��?��CS���b �i�N~q�8�o۪�e�˭-'��� ,9�9�Y�%k����Q�^�N�`���۶cB����ǎhU@��կ^V3I�@�f��]���2�e+Vha ��xh�c�o~���X�Q'�ډ��[��x�>>�pX��Ύ>9�2\t��m7�7�y�x���6�=��p?@�Z���������E�N���3g�9�����ڞP��\Ȯ<Z();w��}�{����<e�� D�+�*��Vȩ�'t��Ff8��o�~G{<�:S3�����[�lA��_�\:�H��8T��5k���s���)ۿ|�`��82S��)��?�*)���N�d��ӏ����W%e0k%1��ΏT	�,w�C@��9K�	1��=��4�}��)��~p�
qN7��B����*��z�ԩS�]]�����CKq�a:o^�.�O���*��ۺu�Nd*���_��5x��U� ����ղ�.���V{�n�d �L:��Obe�pg��2?��;��ͬ-Ro��v����DNSP�1�S��a`ltX�ҏ�'8�Ɇ�K �1y饟@���g��v|R>x��V��kf�z��`,'����XT=m�;�����[���T¬�>�ϟנ�m�(wKaQ���ޮ����<�ڕ���p�W=Ϟ�Ae���yh�*=e�ąv��yF�2�A �D�#=<�������{L3�/%]�,��#��e���{�_In{ä)�@dz��b����uOa7������7VVQ���9,c#�d���*��#�����U��X�L�y�*<|��N��(��͙��A��O�{�\�"Yh�nx��p����4��=f��u꼩ST3�7
�Y�b�Ǝ�x�'ZѮ[� x�)7�c><���@S�Z/������auX"�Wo^��[����R�������ݡ��	���!����?�6h�����<�Y�[�����AJ�XٻiF�f&~���I昰��EQ;
�:��ճ?��T;������|̜��<]*��`g�y,�+�^ ������oɑ37��1v��a���O;�/z2݋��@yD����6�%�˚��$|��!���ʸA�Q�LVc1����&g�wtN����$/�S�t+�&\�k6h���*#rRi����J���8�,j#k�>}
�>�i	F�yB��%���G2ٔ�<u\�6k�e���i�Ih��,�@�P�/�*+Q��S��tH� 
'���K7�2py��P�\���CM�ls���9��mܸVOջq�&��zxW�^SʅA���A=d�[��S��`�-��cj�.`���[[��@\V.[��T/]j�����0Ŵ�տ��n�|�0��h(�{JL�0m*�����P8a�oܺ�����Z�|������dw���>ؿGvV>�>��T�Aێ�R( ��,����r��u�r�*�8��;�����	���|���ADX9h��̞3]6�[-���we��[Ι)�,��	��w���<
�HQL���c-�� 55Ks����Y�Y��'�qձM�b� 5Kv^W���I*Hׯ_/_���r��Yy��Tl�|��������YU�p���u�`�9sg�e2�?��e���Y�Zb�ܙ
ԓǏ�e�-�����aBZ%���X��ۗ�����̼%�o�z5*�~��3𜖲�IRYӣ+��Y�ɋɕ�וm��kߐ�J9��樹i�J:}X�d<���!�<y��O���\���Z5�ƾ'HK�B�ˍ7k���ŪeKefs�ik�%���(37C���1�p�.�^+ϕ�͓��q����+�ь���pC�k�]�P8g�`��`�>��<�c�t޼���[�HuY��l�U�GL�D*�6�c��=���|N6F6��0<�V;�V͕��|Vk�8 �U�+�� �B\�۶mS�E�x�b�i2{0��3gjUg�j��4; r������\���Y0~����7���q,�K������Qj��0i�p4N���sa��	���O�eKf�¹�x�6��m�vwu�j]%DEy���X�y��i�j+�c,!x��/�gԴ4��z�={��B�/^RsG��ѡZ������3�~V#��~W�\%�pȴ��x	�?��?�������_~���Z��� s�dֺ�S䩧wʋ�����X�D����M-��a"�O�TK�\>{RVm�"�V.����Ϙ��Q?��޿�=�Da��2�T<��V��퐇6���S�����������Me��Bݏ&�$�A�:c#�p�k@�\Qd6����L�ʒ�Xt�˝��\^Wh�' B��v�4Ή�] }�Ӵ,�|V�~	��`߼y[���Zؽ��o�Q��u~Q�Q;�Z�ʩ��SB��k���|֤Iu��;WY���M����E1�7���Qh�~�/����)f@�i\�C��khz(�zu ���Fܗ¬�̅8��X0k���3 =~�~��;o�+O?��^��/e߾��}M*+�5��� ���Ď��R�N�������9���㢛l��d���n�zy�׿���I��i�L,��I���4��.�To���D��[`@���<۶������c��L� ��I�J�k����-<�Ա�2��N�!��Vz���	\�՛3l��!d�_O��Y��!c ���h�&pxs���эk7�\F⹺�zH���>����,'9q�\�~S�'�&�k1p�7�˓O���|��G2���Uٷ�=�Gb|��P3�UJS�f�:Y�z��>sR._<&�)�oQU`�6c����F���.�1�E�<�]�KW������V׫���C�u�t<�=�T�Ν�s.PM�c�Jb��k
�'��>Hz�4o�V���?�+ׯ���ɍ����l��.���2�?���,��SOh�_|�E��;Z��붔B�`�>�ltA��XX�P�`�Y���Z���լ��0Xs���0.��s`�t�$��b�X�Ga�-����<��U��v�\�TU.?���$�Q�U��^�F�ǈxu�cBC�܁!)k�@��ժ�X�Iώ��19��427F3J3H��ǔ�=(�Ϝ9��Aa�� ��Z�=���S��O7���C�0sL��X���y�=۷n� �Pv|�G���J?j��g����t�^����$����l��G&�fS��g�q�)%�.��%���J���W+�,^�{�\��[��A](]Ъ}C}2o�"=��E��|�YOd�e�Χ�y��~W|l4!����2 Ǘr�It�${���M@}��/�ح`��[f#8����)�d�C�!�T�-�-�ˋfHoW�m�fCN?*KVm�c�@�>	�3$i��r9�]�c�'����h!���7����[�ƕ�RW��8�l�p�p{C� rg�a�05��$Ro�M�-[!kW���헤�Qe�D0K�����j��`+N8��SUz{�5��z�A���	��ߏ�@8+C �:���5+��P�kW�ܙ����z��������"5\�4�'btlX�l٤�g`�_O�Y�z����x�U�w���2�e!LiX.�;�W
V^�&���Tz =�1/�������~�|xDZ/����<��4�E{����+uq�����������W^Q��A��;g�,'�	��;.@�����?�O~�Y�f�n4OfT�U�w��B3zύ)�]�n4J
ښ�446(8��s�Γ>:���_�D�΂��KJG���/��Sg�O��$h�����n�J%���*e��&����R�Z��g�pC�Wo��AV ��Q��cHʫ�lܼ�s��i܇>D �i�u���ZQ	7�Bf��$+q�h�!��Yx�Cfc���8����L�2YY���Y��0*O�����ܗk�:w����Y�J���rL����j	�\_�Sr���Z63{^��>w	��M�7oި&���C��z��'tw�0*u��;������Cr��yY�n�TW��M�tA9{���,@dYم��G�m߾}���b�\��}�/��'(X��ki�f�b����ߪ�?�zQ��e�bX��Y�k�ya�ǜ3eJ�t��`��+g[˼%z�٩SץK?J���|qoa����DЯ��E9;#����k6I|�[.�=!�E=|��q2�Φ�(���*�P�PH�� �$�6UW?I;La��h*+��G�y��\h&(�*���X�u���~�3�
$ขɠ�lj�y���s�,��q�����8������?^�b���dep�/�?'.^�Lw/�>	���niiV�̖N����;�i�ݴ����>�%M��,����,\Z�%+�!t��	-f??:��S!��
�^cbT����ΝՒe�dX��mø�g��K����l�������e��i�߼��'��%G�={���e���	��0��J_��Q����X����h����q��
���
���!8����94\:���)�3���F�X�� �I0���elf�t�u�25����^`|Y~*K(�Ӓ�(<��˗��㇡�F��,��#�y��׭[�G��350��#�=��<�{σ�{':@, @���FSՒ-K�c[�؎s=���N��;��{wfss7�ؙ��8.�*E���;�J���^��΋����#���}��9�9���'&֊�0� �T()!���i`�J<���w0{S�yPTP_���NNN�f�c�H���sg?g��[x�
I�. 帥e�v_#��`d��iV��HQa����HDX��<}�\�x��%Ղ�%�����?6m��(�cS*T�~JU0g%'gA*��*�^��شE�nH�>˰`� �m�v�`�޽�H�T0�.�_\���n���,+U�^�~��<h�+~p��b`�Au��V��;wU�4����,�Y���R�S���^6�d9���e<�Nl�¾�%��:��V�����8033�beˊ�1�๡'�J�����+Muu�]��}�yr��%��s������7���O�\����5����[$N1ï�KX@���`�&e�тޘ_H��z�IS�Z�}���O.΅x��������61>i���P|UR�px�Y3A�j��X?~Ҫ+!^�$[Ɇb7Z�&Ƙ*1�#O?sƜ��|h�s�N���3��cB5�w�XJ��e��얙�U5��?t�e�O�)��ƛ_Vs:%]��9�o|��DGg��Q̱���8U�;�t���	=dQ�ڛ�ScS�\�,�K�V�&%�n��kT!
�kū��Ckn~P��YV�	u��}�yz;��/�������0��sE<.%9��Vn���P��P�������?�O���J��O{>��[u�aoƣ\X\�ֶNٞ��CpT�H�,{ftBf��$7-J2�Bep`R�ܴ�g
ւ��Y*@���=$�rrd\O`�jX�@�9����9=��(����W$l!�[�'VB�*.!�N�c�G��uu�1::fm��vXw��ꢕ�t�&��'��i�P�2��W:���ɁN�8&)
,��S3�«?�����U�ٲu��������V��k�z�v����?P�Ԭ�i2/4�/��L�t��ę����j�P$��_��Lě�v�H�>֕L9Oپm�uWW�6�oi5=���G��:Hy�sP�+(n��̅�9���4���C���$�R���'cX�zU�~i� �X��P�J�#�ѵ�ղg��U^=q�>C��;Znb�
�T�_����� ��*�C�M�M��@�j�¢|)ؖ��������g
$ӊ�<�����KTu�s2Sׇ9ӱ���b雅�1'F3�6�М��a\�\�����9'��M[˓b4j����!ج��߫�䱣��,?W��$�;M�~���O?�ؼ�T=�9��296��"�IO?sLMT�ܹ]"1�q�W����{�T(&�h��e�����6��>��k�&_O�T�?T��O���c�M��4+��6����"�mMV&�	�x�]�.�x�F�(a�c���Ȗ����(�N�#��(����!�R��7�7����hK}5��&�>����\����nx�\�xI���ckν=��)�"X�UL��(�$�����7��c��p����YN���uu�#�<4z��
D�V�F������H����07����������1��~�zq����d�`�~/��D
 <Bh�p5iF߈�T�S������RO!��0eOG���{*+)U`bf�_�cow��m��v�کf����S�Nȼ>tkS�4�7������r���z��ګ_�SK�BUX�[�6n���Jբ��R'�Y/++��6#��ޞ*�}��ӯ�n���!՜���*`3��ZI
�}�w�ޗ�� ٹc�E�kjjU��%{�yz�/]��.R-M�һ������J}�j������83�`�bl|�j�'PG�\,��h@pI��-g�ļ�^�����P;� � �Ú�S	{ི/hg�yguS�R�y7a�w���޸1�,@�Z3(�w��0�+N��x���`>C�V������B�VЎ��Ӆ�����J����1�M���|�4��' ]o���؄�L89�x��7C,���m13;g��Bv=l|
4��MK��#N����V�¿�� �p�}���!�U27<���a�R�`h��{Ŷ�!�զ�g�P�N?E�n�X��
��$*2ش�L�_|Ӟ�̌j���
epH�j?��������F�QFN�fc���u��hT��@�T��(K�*%y�%|�#�%ng����C�ol�g�)Ǐ���6���"�������K��}���������6e�PB�$(h*��4�!�UCs�KS��r���fAx?�~>��'����!%B8M�2�epY
.ccb�gg�>S���=<��Q��fۖ�Rv���4��Ӭ���'�4�
�d��0+���b� �e��������1�D�vI��/�,�`���nIV��*�Nd�U�f'UR��J\,����!V�g�zz��(�T7�����.��q21=�'2�b5�w�.���a��i�|��*H\L�a 6���(]�����s=�m�҇���,��/�;���P���͛��3�JC}�����L�UhYJ��n�n�kTl��<�uIO͐��eR\��4xlܼܼuG�VY��Ɯl�{��y�$�A'���4�����J�v� `��m��C��2�=^��yľ64�I�:Ad
�y��b�9-Z'ŇtY�1��X/{�-������}�����^���ZMPU�\S��Y�A��J7��y.6�I��O`
�c#�}���V�bQ�)��4 (���i�RAD�"`�۬���7Cs毳�S�V��#�v]#""�����K���W_W�h�WmjRs���`��K���C�P�z��U�<�f��,�<4��55Q�
G\�p�8
>��+\��� =@���[7���l�oH��ܻ{S1M���}�,�G�v�����R�T	C�v* �TMVe�[�쐣G�Hգj;\gξdvL �V��o���"��@D+^��@���,�t��t�w�frB��]�.y_��>N,DNn���Rm�C��,�amF�3`�ٖ��:�Y���rtq����DJ҆.����r�?i��ڤ��T.����)#���XR���� �)�b�l {H=B��< i���fiQ3���nf�NU,�c�;�TC�0��v:b����ba�v�Mjm��D[��6�z�`T\��u�Q*r�@Ϟ=c$�/|��뼜>yԙ��'����I3��>��������%7Fi0�,�=՘��)z��֍�go��RX_?���Q+.�g���^M�&9~r�j�!�ܣ!`d;b[�{N���}�T�w����p��Pp\n�,!q�
O��X�I�����!b�R�KYsë������>�����w��-�G��۽��>.B���,��a�Kf�o k���e�]k�S-�6>6:ر�
�L��ᱸ�����p��) Q���}�����J��q08�v�jRƜi�b$�xF`��5������uN<�P��� w;7����	�B+?yL��X�w��i+N^����7�YZ\�׾�50)$���jTLF���@j�����z�a�sXd`_��P��gO��@�b7oʳ2�l��C��f���	a#"������������8�Nii�S�mVf��֫i&��s�e�Z:�"�MT�j���r*'��urt��U;��΢B	���x$s�Ӓ��jm�s�z_���H�hk���G�ɘxʙ1_����G5р9OT����~F�XW�ͥ''��z�$�������Ң���dY9r���[�4&oذ�#����|���&�v�%o��8�jXb����=�!%��,�/d��iǬ����k<�k�9,6Z(5)�6��Q�z�V�5��<�|��5q<w���_�)��m�M��ٙy���D�P���1ņ� �g�:��s��׾�ا��8�]����lU��h2po��KE�#1Pie���逸Oii�ӜT�ܭ��/+Cr��B��Z53F�q��.u��ԅ��)r������G�̽�	�����e�Kl6��A8:C��P7)Q၊��lD/�ވ����w���V�0hHO��y~p����XJ�*B��~��c�
y���� �m۶��=��o�N���c2��p����ޛ��;_�S6���<�V�?��_��A��v>��%=��/A(����ʧ�jJ���l��6�qK�Q�6Η8�ܬi:2�xFhT�.�s��PE����85-C�Ɛ�L��zESs�qnKw�������� SƆ%/'ע��#�ҩ�P�s��nB7nݖϿ�l�Q���Y�Q�>r܄ME�?�y�&�Y�,t�W��V�R�j�i�Б��Q�=�zF�qJ5/����6���2
���d�*�_��7�EH��8ʇگ?�F}���m^h�:W�{F(B�,{Y�[{[�\�vUv����>�F!���_�k�U�&d����ߐ(��Fr��W�3��!�������6��=x�)gr�YA]�=�<�D�ҍ_
����@q\���յ�+�5�d/gX5�������@��A%�"H�8�gh*�<Z��au�99��f^�y�mSݯ��-
L��}��3"����&&�R�|��uk������X2>-85���?�v�?��?K�o��:~��Z��� mIY�5S  q�I�����;~Ć?��8 ����2;4<V^���a���:$6tp��)�Q6�6�B`�{* �Q�G��!�Ox&Q���������=O�?gdp����R��KLl�u]/��DM�0�PŲ�6"�:o���M��I��e/�N�:�*8�_�Xh��%�:֜� Ȃ���r�"O,�Z��?�T���b}:�Mp�aq�:r 3����Є�W�b�F�
u�à��.��W������OZz���޷l٦B�AOH�M�@0)wƻ$7F�.*J^�̆zu�{%%5A�"C���L7�SOn�EKq�ʩ���eA�ǝ�j^��;�]u�7���R	�Tl�߄3W���L#��F���ڰ&����δ�I�i2:�� �L��/�����Q#Q|G�3��
��	�����RW�U��>Ňajz��3V|S�P��cپe�b�i�u�VC�ٻ]�ِ�=0���'O�֎V,Zl������7nUşT�b�yk@��mcd��E��
�!Rxz�r�sMI� h��i!#{�f#����746F�q�g
�^l>99���(���ZDͫ���%+Av8q���lEkѺ8���f�9ry�Y �9�����xhN	M���dN�C�z�h�i�hq��媭����KbT�Ғ�u��-�[�%���j���eZOnfZ���=~�%����mN.���}x�ٳ��=RS]��*e�6����˪$9�G1�!;\��m
�We��"�N�R�Zg@��K;��`6�4�{,��A����J�۔%���Q�쁕���.I�q&($�s�6[ܮA�驹E���^Y��&ʿ�կ˃��m��|�MsB����Yh��1x`�1N����a���3]��E4�z���}rilƣ
������N���t����o����j}T^����y|�S���a��z���-���6��$p�.:���`s�|�%��&y?�ƃ��V(�����^��Ʋ��A�d�����>u�~;�����H_�\��.}aZikQݭ8b�<�u$H���P��ܺ\��IyE�>�� ����
�<�����f�՞�.�Sa�)xfzA�V��_Ń��U��Ip��.z�01ff
N�$)ض�>��k�&�1�J��8��SM�Ei�}d�&35ٺwn߾/�)��6ԶI��ꐈh����ޡN������E�P�����J�5�y�j���b-9��;a͌�0a��C�}N�J_�V��������A�CxǼ����1ﶖ�-*`����]�R/g���O��.�E}��a�l�F�M��^�a�1hT*��iw�͉�9{
�i.u]v랅�ʒ���a���`I).ޢ"���  '/33��F{k���޷)�r�t�e�K�ñI��oHL���j�f��iLx��|K�c]�UI�H�Y��O~�+��z�x�7 TZ�;��٩�䞩ô��
�-P[��4@lT�
׼�F��Y9�����JU�}��3E�
��ާ&��/6��p�xW$ۛ�jl���������XP�vT�<����={�ڄZ����6��ד�m�{8r����Q�,��:7{�1b)�fY?�CNM�Z��u&�@�R*m�z�)Z$��`��B?:��!ƶcu�8ak��}D���U�ÿ�L��;п�,:*Ii���T���B~х�c:k�邶�kj�ٔE�b��-a�P��q�Sy�7!?`�`{�C]�$���e`5;8ԥ%����A�mb'〺�[�檶�k��g�>a^3�;T :�Cܶ�H���\�vO�Z�͛d:��^�W��W>��Փ^����_��K���-e�*�cr��)��UQQ��oB~؈eoݾnxtx̪3&�G*�&�0N�"��3D5�z��r-���/).3�H�޽=C�9w����iŗ7�\��.�s�� A���/�|��j�j�l��ajG&�AE��2N��"0�&!�Ev�M~��w�@d����(;y&�G,���uR�eD�R3��V��[�d�.Ft�(��1�S�w�t���᠌�Y^2M?=7�3����D��Y�_���\%�a�EPZ��KV�]�`=צ���Bs���>N=��U�z$�V.{0��fY��UՇ�ɱ�o0�R)�����ISÕ+�ʭ�7�����YF�=��K�v��#�9p��m	�����s���\ܱZ"B�K����AFGf$7g�̪&az�����Fݱ�TDǄ�k��j��S�z��d����~p�؞���$��Ԥ[�#5����Č����D*.��߯�ҡ�d�r��.��O�:)L���eppL:.G��?�`���g�<�䔕��H�qw�7�fJWG�	&���ޱ��uJ��a�bSd��p����`���y�.�,cm�O,��
�d��׽����gF����U+x./�>Q��g�W�V7^a�Nk��`��uB0����[g�����ͨpT*����7h�b�z��{�9����˲

j�;��R�w��Q)Q�sz��I�fyX^���8��b��Wo����F���@q���b�w�L�:�Z�ܢ����erb�4넞��=sL����bٽE;�����O��X�+����B�K+tѧ��6�GK��O�o�d8�xŋo~�-��\RZ%���ln��c�iji�U�e	��
���o���Yfv��}��cvY;	F����HFZ��h��{��m:����P����|�8��J�)��А���1�^-�,�Ɯ�ҩ��p�N�6r���x��.e�X�@���=��s��AO�ŕE5?�!Ak#;��L'py\����{��g�M�{4�D��&*�U�H�[�t��T^;~�0�
�_|Y���~	�-u񝝽V��J��M���t��I�*P�U����8���C�� �V<t�O��IJB�ܸ~�rh9�@�w5�v����Q��IOI��jhj�r��������+4^X5��O�E��d@	M���T�d�!=�|�����I�T�[��v540,{v�SO�HJ�������^�'w��G'GM��,�j�5!A���2���?�������ֽv�aN��I�Qb%K�<���}q�\�h�o!��7N�{e��~zm�����Ĝ�k��Z�����;��(�X���#kS�]���#dļ,%N�!������Z/`zV��OqY�C�
�$���\\|ג�t�lHH�ʲZ51C6c��p��G��q����b�ȼՈ�X�]�Խ�wԋK����&�^�٩'2\>������á��*y n�餿�	u���dڳ667�g��d��K��ҩ)��9r��i�Y�}�X���ʦ��ҤNU��i����IIy��רr�V,��;�Y���/ݦ޾N�PE��رI�iu�;���nl��`�O��¼Z}�z�[��u�,��hi��E*SkC:��-gV"�0���K����"
�wm�:��o~~s+��fP�������
���q-;e2�`y�M���y�n>�e��˘j�$W�H�z�Ƒp��$�����
��M,{�-�����3!,�_*mͽ��c�-��,V�T��+P�(��4�sϜ�ώ�[�n*�됄�G��^��v�����\#���ge�J�~V_o�t*@wI]S��TV��#{�Cd1��P{&N�����Vq'7n�W��h%�a+S���X�{P���7뇕����9Yyr��M+m~��/Z��������ɡûU��
�j:�+����بH��=|��4��G@�w��]+NMM�*Y�4C��Q�b`��,<������8�\�9<��s��b8������;�5�0��p�HU�>����M���~^�p듬\��J=�	w)'�k8�q`¦�ب���=c�ihe\	�B^�K�\@5I��ȰzkS���2$�����TlUutd�͡R�CL'##]N�8e!�{
�����ܻ�����cD���Ⱦb�������/K�: �M��h;|������f��_��
}����\rR6lD�j6��U5��������B��6��;*?��3�ǃ���Cd�m�S-աۨ�X?u�p���یp���ɘy�Ąx�ԃDF#**W�|��:��5r�݂K���A�3l�ߌg~My�8�P�����I3�����7N�����I��0;��0Gs'!�X�P��u/j=�0�xy�fF���y�������;�|�x+gS�uJb���bt#�:��[z�>�!Ȓ<����W^zYq̤�W\2����_��nL���K��qZ{��F#�u���Y�X}��QQ!jf�m �}�$<,J�K�ʹ���뒐�$��k��R\�(H[q��8��ɵ�er|�X����$3c�Z�:7��˲w�.		0MD_����jB����v_/������(��sg��DGȝ�7��ED�&à<<@�[ne(�yN4UcS�A sd:dCr�iC���S�h4�*�.W��I��!�hv�@�u��⽎09���^�y���g������n�*j1��]@�.[�~[c���t��iC�����,]LN*������\�I��׮^7����>gy��]�89t��.x�.�5�h�l`���)+}h#x7oΖ��J��o�ݜ��z��V�y��Usn��a�!HD6f3�2N��'���£��Q�<n���9��)]=�Ɯ�p��)3MS>�Ve@W�Ⴧ,����^��d㨮X^���~���P_�H���%\�kzb^�j���Y�B���}uM�u$�������}+.��"�g��sP��T{9�L�&�֖�r��I�,?w�#�;��m�5���u��z`Q��7`b���'c
��i�n��ɵ�z�r����ܓ�s�sY%pյ�ˋsh���Q�Vi���,�}��=�F�~�2qy�|�ӎ�iP��lS��by9T3�T��̤ʁ���sgN[����͙�nq7�����1�\���@��G����fuO�:fZ�EA��ܲ���)$�tP��o���T!�ХZ�@��i�h���f����P�"q>95o�<��8@����jٸ1]?sm���	zFj�
n��նH�:�*DM�-�����:%�)�Ⱥ2w���F�ojj�
r�E�[��Y(�iTt��;�c�+C������	��Z���{.��K�������-�s�*�K5��,��(X>�K�6�!���6�r&Hh����4Ϛy��
_�7C�x�W���M~�w��{ߒ,�R�)yTUc�9����^U��MDX������
e<�qa� z��uijl���Xc��H��W��sE�8`#HH,���w��頡��&
6���WM�e�,{�������b+�Q\e���]8.>�ʥkUHvV�=|@�zz��Vύ
�S�)��Xo��'��җʇ�2<�ok879#e��ef���Y��^�]5��׊�y�Ν3煱v�j��~)(ܥ&,��(��h�a�k7��3V˶(?���U�9&�o\�*Zl�@�1�8G==Sz��+65ֆ���c�
��ʨ,`2���(\E������䔎~�2YjW #@ܿ3�Fb����&�ka���T�뜐����j�H�k�+��G�j!0��{�ژJj��9ڔ�g���fu�~t��Q��s��O�?e�):[�<�EVuG�׃`ce��p0II�r��A3�,&ܞyz�A�r��}K����׭�	��g=vȞ��i��nG���`"�yx(�"��\/�c�*�L�����u9r�ezzdb|Z�b�?m����J���4��0e�Y�[��[�B��٫�H����J��0���{��q�~�0���-���8��Wg �����w��n�No�3���f��o�Rr��������.�{-y,<Y�T����u�;�"�)��]a��`*wL��NN�ߐ��Aڑ|#ZS��t��܍&@?��?�Q=��;!d�)	�J�Sw������=
�=�&�ώ�9h<uM
bW��ge��͖k;�����Mt)�3ǢSgD��o~d�ɱ���u�����i��FԘiy}׈�z��9	P���jʘ���̸����d���6ַX��G=Ӊ�9=���/\��^�QLKߠ���BF�����Z����;�ٻw�I���}l6O{g����m���W��6ȩ������6ZH<�v&�38$ {��˜ ����0�����1o.H��KK&L�#������x{��'k�%��[fo�XY�S��u���~7�z.����{8@���t�Z�)��b=lyE�����A��`aqF5�3���Njj�o/���XyXYk�F�IS�CP0Z[�(jn�C������G��R�H����V�6l�g�=c��^�a�^��Ss�e3��}�W_�v���+��ݔa����L�&�|76:N�CB%@�����+c�S�qp�K��I�:9��������[ZSy�yKR��Cz�,@�e^1ߕ�7T�w;��ަ͹~L|�4��$̱��b�>о���z��p5�p}��	��^-��k�_l���AӭE�:c��rq���8H8�g?-�J���⪾�����e��U�F\�"˽��x��=׾�A37q�&� >�辴��ø)�Ѽ���`��I[����֭;� /��y�R�O?6@Lu�Ǌ�+N!�G��X�)�W`vnQ����$<4J���[Y��_zU7l`����c�v�r�3F���R�&��Ǫ��ͯ�,�y��S��kO�%�����ZĚ[ddtLRӒ%sc��w�'wO�T���]P������n���zJ}[�L�e��!�6���w���TMD���m��Ϝ�,ŝ��F{	��V�ЈH�X�'��0u��wޓ?���,M�ƙ.�K�6}��B4?�=C0���)���o�	�G����k���4��*�sO,�pGǇ�'mC���Q���lj���ZX�h��n��R;zj"�ͣ!��`��S��5�+�Qf�͌�P����m�8z��\�芙կ|�������{�K<��Y��UO!������;
�[�3�n���k+���D��o�LS����놂� 9}�y�W�_1�My����)�&�1�֘��'J��GD�^��ۖ�ƬS% s��pF��~��k�Փ������1[�j���M
w�Ilb���+Vk���׊�~�_X�=�s�@��-,;������9ռ}V]����}��� !>ƚp��ض5O�V&Y�֋��$3KF�D���j)H]h6�.���i*�7�nq��Zc�[��V�>9�D�Z]]�
	���v��s*T6:l=eC.��%* s�S��ϑ�!�!�`�l��
[7����.IH��)�,3,�ܙW�5����my�dcf�e����$��HmC����'�"�M�o5�/��Y�����e�����/�ݏ���+2��|Ѷ�@��l��{��@xHRj�͉^Y��ڮԔxk[���Q�}���-�K���>z�Z��u��âͬa���Ԍ��F���.�u\�Y*�-].s�c2<�h+ƦF���5[�e�-��o�^��hQ��N�����]�~�����}V�ME+�Om��`����mpU���9u����Y�q��-�eи��ҭ>iS[����̇�	�.)�4��m���:&&�0(#�N�TR�䨨��@�V=�7$x4*�0����������ܤ��pcY�D��@��Zjnn�L%���4~����bPzÀW]Wm������Sj�JH���Ӟߥn��u���}����Sa�"�5R���x��f���|yTUii�<�&����7�)�m��ɮ�Vc���N���	�������t}c�K�j
�:{���j�`�j���B�աa1�7N�w�x�ƴ�/����3��Fs��!�(�`�W�kxP1*Igj�e��(!�W��f� �P�������FuC<n|̨U5�>²<�f��g���4� �����.�{�|�>����3��H�[֌����$����^	�	�.�Gp���=g���Y��b�P&�X�S�����s�9B賎�x�V�7��=
���Ύu`���.U���m����S���.Y�i�] :���lݜgC�jjJUK�D�Dʫ/���@����t.��|�v1��*�!/�.]V!��	`;�v��������:,�>Y5�5��_��쭺�u29�)�
�Cj&ib|TR�l�W�
�Z�	)VYUUm�HB\��K�z���@t�0���}���LH���ݻ�����q	�)�6�r�p�GGG��Z/=���e��ֆLe��ҫ��Xs/E�~Ϟ}��w3yk���",��P^<v7d��ͥ����{�bi^�&��7��}<I�TK�$�&+t����M�\R/S���Ç)E��v���o���\�!� n��m�@��X5)ĥ '�PA�;�p�3s�)O?s�Nǃ{�̳av!����"'*CO��������w�p�#�oU�3�?%;vK�
c���X��W���d�맶M��mڔ%�^��''g%ZM_�:?��U*��Fʨn<x˼܄h�[__�����@9a�٢f���=�0�GZ]]e��	q�i��Y��op@i^=�!�oDs�:M_ a����3بBA6����i�c׮]���6���Wե.��8���k��q�8�0ߨ��n��^^�sZ�T!����Yn4yG�1���ȨAńO���Ű���PT�[�@?!�^�	�3���&�M����̉�����a��`��K:�?�"@8%�I�)�9[�CKJ� u�5�� bq������:�t����I�2o�RiZ�YH�
l��}&�T<ܹuM��@�L�	hDrb�x��ʏ~�+
�ԓ�=`�[Z�2@~|�1��F%�dYy�v��_���[��c�y4j
󁖌�U�WzWπ=�ᢝ�v�ү��07*i�	�r"�~��5�޴I=�g���!�;��-j�X7f,B���3uL��uG��)7���QoF��T����+�g��U�*^���2��a�t7;�7Be|�k������	s�TPaʆU���g.*"��D������0�.�� ���Ǵ���y�FI�bF��f�ٜ����%�b�*X���YD�֐*��]������0%����)HG��W���uf6�Y�k�zX��9��Y����oZlqq�b	O9v����B����ԉ��TܹuW*V��ؘ�+7o=Ҁ
Szz����ʐj���e�?���n���n0�����ꢴ�5JO7�Ì1^���Z����&<_Oo�i�J�vh�)}���~4
L/:�--MVE?DeE��~���C�Jp�;O�
X4�뽻Aj���cq�v;���'a�y�i�G�\fƹ�y[[�>48���ň�!q�����B����a��<1aus���2YT������_��,�t<E�����;T���>c<�|-��T#�����P̙?P!�lc�Q��5��Le�*t�`��Y?1���u�WIS$%ś�s�ʧ���U��1U��>�f���g�0Kh��Ҙe�~�o-����V���>s7m�c�l��Ze|�W��)I
�������ۺ,-���7#�@lU�F �Rl7(YST{Ęg7�?d���9���'W��OI܆D�
u����"�z��>Єs�,j`�JՓ	���ʝ;��CA�����F�L��C�C�� �'B=C0��Ҋ	5��5&]���	J�ڔ��U��ppp�RdT����,G�y�NLM.'��y߾u˪ W��C��_����A��w5�ME�
͂��m*�~�M���� ^�W�(q�z+ay��g����Ư��?v�y~��?��=0�`�
�/^�T7���J��s�������g� ]�z�W�A'��i��S�Y��t}�c�u�5V�����gtH�	�#�G�?'�	HI�W��/�#��*��"�����Qo�۷�˦�;gk�bDʉὢ�ן�LsS�<(/W|e�E�.��ZZڬ��C�s�)�a�BE+>��3����R_�<���1�X�!�L�-��0��cYX��Ӟ����PGc�ٵ�.my��g�|g֦�"6�*&&����'lnj	b��W����G��#��VOx3�Uh�
���1��#�95>L��+��9�����I1�ssKzz���TL�
�Dr5��`���Z��h�C�e�b�!��/|,�]�&|Y�FOgs���G�V�/o��m;"o��7�����q���N;|�.I[lL��4u��<G���g�?����S͔��N���¢�W��v��Hգr����󍣪�䎨��L}�.5Q�?�!S�	i�OMJ�~�w~�+KC�m�6mC��w�= 9�y�7��o����m���MC�6���5��>�p
3�ӆ��H���h4K�������M��\Qo�t!Z<��ĝ�:w5� ��p��[�5�Q��ߓSLRӋƂBӨ��)�?-## $(�p|��A�b�31VP`�|e�Ţ�"�3���;��4�(��bբ�		S27��_A�u�F�Hp��h*^ς |���׫1b�Stڀ��|���v�H�4R���my0Z��^��������!C��Z[��S��X���f�,��C��˔�7.�@����lx8��GdCr�����>0�/��1Y����>	����|�z{x���f��
�B�:���}ϸ�!uv���[ ���G����9-�B>2܊&_6�gt�!ƐvLhww�	�޽��������L� -��+{�4Q�[[�­<����8���Q~�������k�~|�c@({�70"��h_�����cc�u��`y��v��-�m Η.�� 7@���zR�'N�S����ukr�-Q�ܐ�Q��x������	�r��!��՝FNƁ@�j�����yX���o���	�뷬W�$6���f������a��s�pkVVU�`�����`c�}zQ�z��p�v�<�|S]{��!ټ%�:�.�!HIMR�n�ͬWO0I�UA�]Vr��r�$�����ژ<O�'1|`����a�5|�Lꡱi��˗G�T�_qWTD��f���a��  ִ������6&6�bh5�uf�4���*�vY������1X�uG{Qـ&c��|�-�WSTi$$%��c:y�����5��x�4��-^������x�W_�#X���l6M����ŋ�����%��%�-X�[]�܀[i�àu�<��q�kj��6^q�c���X6*:_}�U�K�q�	t\�ܹy�L'��wh�{LS������259{����r��E݀z��+��`#�\�D2UX6�締�猑�_M9x��Z�t��*RY��\L�=&&Yr6剿>o��J�zG��a��䴾�uR�ਕHVP�*!���Т�lc��*&c�0B�0���U-�?^,�3Jw8�L�ݱ���C�Bwh�q3�Avg�1D��WO�Ѵ-\�?>�L�Ԟ���2�蓈X4~L!RR�E����fB�(X����{�u��m��w�Іf��9��!KV>���^�U���4&�D�Z�*3	֧��Bҥ�!F2�Ee#�	D�C�%Jo�����WL+���+f
	Alޔk����l�^Pn�F�U/��_��8�ɻ���xo�]���go�y���F�a����5;�$�<�����֨# ?���}κ��X_��M�:B�O���E5pFP��EZ;Z͜ӊ���
"-�d�"cg)�ڷ������v�9��L���Ԯu)�y���֭&@D��g� �w�,���I=<6,'�:e��H���!cV��´���0��ڵ�VF�pt��L	��nZ�<'7�,���[��Z1�DH�X]]zr+�/pjIE�M���LqX�nh����z�n]���F��`�:=ynI��B�I> i,��L�mp: ��f�!^W�B�{�#����ޱ�(��a	�G�h;��>��׬��DK9�{
�tfnZ���-�U>�|Y��&3����+V�N�u��M����6U��z"�2s�H�jY�qDt�Q{��s3�i`dXr	0�A� ��<��lLۨ[&��o�ڹK_�Ÿ��zLk۰tJg��Oꆤ(LIOQ��uz���A�)մt��p��a�߼a����w�j`�s{Sq�M�r0�[��@�>�̈́��s����iCfG:�x��!4.S�O������c�uxT�4�6�g���9v-l����`�BN���.3n�JzY��G��n���R�>>~,��yUΔH��y6���QJ:��"u�v�N�[�u�>�%�
Nwl�&/�=�.z��ߓ7��E`ƪ��4ɑC��H�ae�L��(�Q|������y$|��0c^���#��}���I��ĩg$$"^:{���	��O��u��a�ғ��C#c�V��z�ݥ���gJ#04�6�*O]�VH�P��^PXda*Ƙܡ�g\�ujv��U�eZ7�^�=3��UQ�\�d�� � x���Th���
��#HV�l���Ҍ�����Ѩ|��v#�p�����P�E���ۂǿ��-1�!��u���^L��rJ'88|ai�CT�Y��:�-��[�-�����;\�jŉ	�u�m�7�f�c k)	U�̬����M6L�FF��]�1�}�0)vxg�nܲ�c�[sJJ���׾�		So�=#�}�WdJ7���F�j�U��Y����L2� I������/�yW�N)2�˴�̠`	Ro	/m`6�3́���&6���>�,g����̫m�[�}Vn}�R��ћsP	A�'DIvN�L�a�\hlT����A��-����F��	�v��ޱ�e����"��B����qB��u'&Ƽ¿�˿����S��g=V��˞�l޺M�6�Y5Nwkb���	jnTS 7n�K���ʼ�,?Q�施}B$$2V�*�<v��?|Hn]�D������~�Yu�}��\�H/-U�}�"(�%v�`p�c|�ئe��V�\`Q�N��GZ�ر�r��U�SER�D�S&|0����/��546���,%��\�_&���2;���W�RZ��ڲ�	������,�96e�(yIi�j�m
��G�ڢ�[��S��鐮�ǎ��?*K��6=�t]?n�3r��Y�ȑA�Qz�[[��l�ݶFP��2��
}T�.�>��
����lW�Ta.���//I8�����[- S�Hc�ضU6*�#WZ��i}��j�^NiL.hR��_�w5w��p�#��V��G���(��k�gd�_@���I�z���U�K�cYMdF�LL�Դ<�����eϠ'�BZ%<�K��[�j�����k�� Փ�����$/!iU ��"����z9�N�q�,'VO��3;7GB�C�a�On/-����t̕������$�i�P����J�Z��ΟW�.����'���0>wr�f��h~�'ޭ9zPZf?3� ��m��{�Eg��MS�Fm��1ိ��%^7��q������#o��i�������+����QoÉ���NC�inֈRhX�j���;�[	
�JSc�z���2�Q�B�4&�)�D�p�8B��k׮���$��!nۼ�
�f:\r���������ێ����_�gd|dЪE�3�Hefn�2��S����<Ã]}C���/4�xy?���`9��I���=��H=�M��m�1#݄'Dm7խD�qM�N�2OM:9k��ƦzK� \�vU�C���9�%�O$�����y/�kl:���g�Y��(�����m�2�b�Ғ�i]�"#�쏫p�qF�޾#�U���l�Rs�����d���n�X3*��㣒e�K�
LWg����U��w	�_�z�Qz<+��:�<�ёq�z`��s������Z��>�(m�]���%Z���������p̒˙�s_�r��`2����oL�
Lp-4�3��ﮠr� ;�K�?��&�||��v����Q�i�]��C#�E13��������{e��3H��{e��Ʌ~�Я�zx���?j�S���*�Ք����_%59E�*���4-�V[^�ﵦG�kVlc�ϑx�7N	�ƕ^Xvc"<�L�a���T5��$`�|#�C<��YHz��7�|�����~ʮ���`%=_��[Z�k=.>��c�C���`^'�x7D�-��4��8�`|R�{{,�����~����cq�+F�
\�fd!f�>��󈈓�0~�4Ͳ�h�{�T;������,�O|D���� n�R�Nxv����m�ڸIj�_������n3�q"�'����`uw�j�!��b�S(HT�=e���&9w�f�K���)�S�9TXV��(X^�ۀ ����a�Гr��}y��%Y�+�&a��(��ri�7�l�CF[�>U<iz� �,:_?��vǎ0NBH`��>@515�H;V�ɼ|���װ8�-��]S\FM���>�,�;-T��o����t��a��U�1��Qxd�3�O�&%�Q��6�~Z�VKL����2�Щ����`}]mm����j��<����L)�Y�0+����Q�Ya�ǰ�xz8��k$�3�����,d�W����s \����fB˹�
�۝�����6Y�G؆�� oS�H��
�͛���k@��Y �BC�ъ/����_~I��S���b��n���8���Y���%W����������Q����sX!Ϟ>%�N=-�����6��h�U]�?���iH5�g  4�",��Y�t�����8Q����C��o�X���Е�//+1��w&`���E��L��[oYk9��i��^���q���e��B�����,� ��|�uX�����8�����9<��N,Ӎ�����h!�i_Ô�����:|��y�l��{6�WRl��uYh�YS����޻V�hp���M��B	���Ojq,"�d2��<���A�;�_5���}h��6o�I_������s��=�?�c�ėU���,��>�鱸���d�ŗ��:p
��˲
YEU�?�[��n�t-��&�������#+B��q�c�z��u�����������`�rr��l<ͦ�ow�Y@�B���d4|��&ttK�-�������S����駟�������k{U+M9��z=��C��Ɛǉ�EƋ�sm̉F����la�^T��x�3�Q�����ܭ�cR7���ބ�0���2F]�
��\�����_��V����4�n�A=��?��K��t"L��J���p��o����F���f�]�5:t�l��b���[��o
"_�қ��9K�_/���Z�[
���������'G�WV�zxy0���a"&v�\�����,�sP>9���gsy������&R/����E(x@3�ã�Pˀm�� �����p��b� �i�`�8z�2���Et��$�|����PFВy�x�}�9(�3^v�t�:)t6cV�#��豓���i�س�U���R��l4�n?X�U����b�0W��ܞ��s�f�����2ߣ}�uĴs ����|#|h)�5`�!k�6b}�<�����m����ޏ���Y?֙{
�� ySD\�B����
)�F'%.6Z>>w^2�6ʮ��,�PZ� ���A�6I�SO��ד�fV����0F\oc�[U�965+/_����kRQδ�~IMI����o��hY׎� ��I6h�b�M-M��QϜL��֪ X�8��Pa����^�h�v�mD�z/��As~��[V��PWoj[�ZR�������~�sFG�L߈�m�7�811/���0y+�_���˯�ܡy�?'E��D�\|��7%.!��8�ϟ��}�`;8��#B�otB��yf
�4ʆ��n+����@�d<���ўh,w���wG�f?�я�3���/V!�G�8�\��X\X��Y�L0o��Ot� ::�����W_���,\�_#�Ju�$9>�H����<�

?���x��[ȁ��^����$).)��v��CG����E�!�u)���iq��eS̬�$� �@� (��L焹�1���zT�;Z��j�'���rN�:%���E+����ɚ,Ξ=+w�߳�FZ�^��vJv�	=n�� �L�S�=�͍������C�yIJ˰R9�iQ�X64���E=�7b�?������wX����N�o�a�n�C�����4�aM�S�\)�ɆI�
��}����~�����U�)"xn�B���4��������C�9k��q0�z� =�}��!��Ξ��P�)"�V���{�[�xA�.��_��˥�{D�cm��91��+��R���Zr�e�!�D*�C}]r��-���^���ͪ*�%J�L��6m庹�k-RJe$�1�p�QU�8���奦��`'�;-����$���L=������dsӇՔ���3ϮO�>&:V=��5w[M����̃��H��6��j
2�pմ�$R\Z!5�1i/���`��'/=�)ycQN��s{m�8!��r�$��ƧJ8�I6\}��m�|�3�yѸ�i6�#�����M�P!�	l�8����t>�3"(��F�;��v�o�\���6�͐��x4?�227�#������s��:�L��7$M����r���L���z؀.*^V=|��䔎`	���È+VV�<�b�X]P��l9q�)��Oh@��ol �l\����Q�l�y9��N������R��hL`q��U���f� �և���C���r�2������J�*�D��z������C�26JFj�X;;Z��;pPZ[�-�t���Z��1�3^u6���󌼆�a��Ǩ�J�1/�018��g@��Eg������;|��!@�d8��z-�"i'�ڇ 1� ���@#��˲��	6BF)�Y���7���{(�,�|�=���U�,,˷��-�Hߨ��!�z�A���-��SO����	�����L�drvA����xyyzy�>�{x����Y5Ii���30D������l}w��Q��(9�X�b�5=�?��F"%�Z������LϰM�� ���A���<\Y�,#��N�x�<�f.���Dh�����7��s�����g�VW��m1��ǃ�K����40�u����($"�ʜ¤4IK�ѳ]�i��]9�&Pu��këB%@1#�o�MZc�FF��}�J N�9�4�@�PrR]F�k�9G�s��L����1�p-�
6����{;����7��pb2�U,N�	_�Up�a|Ʒ��m�ټ�<̆�F�YT�������!��q��_},%�-2>�)��~��c���\�|2x���Z���l�}Yͥ�"}�EW{���w�7�`��#vbF��VXD��d�:,4�͸S��
�睪�.�����4���'��q�S0�B[���ޘeex�A����"��$&%H_�||����͵V116<��: �-����lݬ�*]�u�P�,*��$����i\��� ��1�JL��p���� ���V���H�&hV�k[��,8��3���}���ؔ.��322>�u�cc,���E:��	��ήu���#A�������;dX�%7��F���u>��s*���oY�\YYcP�TRe��ۚ�]*�����bnu�斖U:�H3�*eK��O�L��� �9!Y��'�7>1l�0M���z���)�=��=�;}b�!���"\�@��Z���T�;q┼��{��Ϝ9#;�_�<��)ή�[���PR�0%"���c'=��Y7 ���旬�L�\��҇�1�VQ^n�!���Q���Qՠ;bn��b�{�<�l�5S#r�r���N�ߒ�Q����'������&몆p���3�!���}�
πV�sm�A��mx�x�����ʊ�F�`����.�y��s��|�{�3�E�!F�&!�Vm���ha�n�%a
S?::nk}Y=���hy���!�sR[�&/��
�8��A�Y�V-8�d��㹤�pŝM�=�
 x*B��$E�P�c������bu�PG�)q
�@N��>ћ��F��)���n���h		>r��>U��R^Q*
l�q%����ܮg>wa��);����=(��6�)�\�L=��hF���b/b���S��23���	��l.עOrn~F=�����9\=���ԑ������O7!�m+�7�F;���T��3ʥK�LX�L�5������f��a$��ZyfRB0֗�c""��_~�+E���e+A�ڼ�3�4��>���cq1B=�6�@3�uu�m��h�?��?�؄dy������2��K�O������#�����%B;��l
U�Qͷ���֌��8`B��� U�q��&�g o3*t�~|Y^x���*���a4ά ���īB��*���ü���[-�����J�?$�~zI��_�Y

w���3�}V��&>�3�ʦa��"�I�?�/BLx��f���#��S���Z*7g�	��˷T[�Z75�����O%)%Q�W�b�f�~t��gٺe���G��e0���|L�l��F��5)����T^Z����K-�ES]u���������	zp�T;�h���!JhM�hFڴ������� V��;��D��s�I�|��S��k�3�T��Ĕdy�젣հ^��Uʕ�˙�^�=�I�Ь����ɠ
��hY�`��������Z��A��ʲǓ� ���F�V�{�seU5�E#�To��@�+r��=��
���M
DW����������F�8���O?�b�Ȃ�U�2��:�A2��ǃ5(9A�����ޅU��QQNC%��1���द����@pٝɌ�Vz�+���%�sr6Y��Q��i,-�Z�tI�����v�ٙ}�u�dJ�O����?:]�eL
&�RY`N^���6�-��$%2<ʮ��Y#]�>~>@uK��\��b��j��������G�,�i�f"p}�F߀ 3韜;'?�����~ �������o[��K_��:K���gyP^'��)�p�f�%h`���^&�^����׬xzz�h_�c��b����c�}��Z�/��r���Ŝ��f���KO �F%�1�D�8Uw��9v�j���t���܂�����7�96�}�N��E������6��
�8
�ֶO*�oL��$���LЬ ���O����6r��۲îC����i��g;��А	����a��N�K�]����ݳ�x?9|:���Wviy�15��V�7��6;�Im�|��G�@�~���0���A��(^��d�@L,
ain^Ν�@���c�Η_{U��ۯ��'�32�?d)�wUP�+������W�~*�ղl�Uk\Y�b
�6@(�j�a��z=+����Uoo#_/n��A�TTިM6�R�l%#+��$��-rN�륗ΨW�C*+�mzt�b�i!���"��_�v�kׯ�wץ�e�#���@�b�˦�>x`B�p�3��`q��sF=�`�|��ðq|!���E(a�(��iE�yG �oL�� f.x��e�Ŝ�� '�3Yen3&oR�yV7��l�a��D[O�"ǜ;�*�I�(��::6�fzn�;��dԤ`�3Dt��+4 ��(>�W�a�
�a��P�&&%�s���k���X�bIN=uZ��<�Z�M�L���G������KN�f�r�L.]�%s
��.�0��\^���԰9��V]^l�M���+#��ZU�i�p$�YN��/$�+�ث2��)	���M��,��g�[#@��p�j���G��m�pXx��%|�+�]���_>��kV��vw{Z�����{��u]g��W9thd�@b�b��%�0�d{my�;�g�{���7����ٲlI�D�")�")�"%0�	�@��C��ޜ��{_Uu7��-~`�޻��s���Ө�R΂�ʫ/�� v;�uB�6�C�V��S'��kX4
����v����p�.Z�T4E���;���z�a�����wI�:��f�F��4��c1���]��z��34��eS߃uj��-��-�Z��!��ݏZ��9��x��'Ō�8�[��]��+� �`��_�O~���ҕcl���{���x�����t/[K���XF�����/�+t���O�w~���d��*���j����N�	ߓ8g�X�'p� }�Z�|�a1�%\���c�q"�u�	��[L��Fd�	�W�E�t�O���Ƞ�ēh�n��ʑ��tjd�~���U�x0�4Đp�x�̳O�	@�j+�LG��x$Sɨl�"��TC���A�u����:�3�i�@��ρɂX,S0�A۠��DhK�6�F��2���(
�	߃�-%���BSI�\��Q^�~tʠ�|�h)ӿ����C=+"՟��k�&��� �p��p�"��3��3Y�����c�=��~�>���鳟�_��Whw|��Ͻ ��7�N_�◩���>B��������D�,�ڐ��ܖ^]�E�g,�sLBG��h+��c�ŞWB�j�	X�����ӿ��y�C>�5���[��e����6��D��4�iJE�0����I	���B�3l(�M,�����L(p�;���h���w:�N���ڏɦ�2_/1� �-Zj�bUؕ�*R�7y� T���x�U(�osH�̰���n? 2�*&E.��� l�^Kp�X�P�vz�C�f��C����#����]K��$�4j� ж�B�͎̚s�՚��.�%�����6�7
Ɲ;＝���/Ig4x���b�"�o��K���k_�����w�m��]J�lMjz�O�T���P�AE��2�-�S�����2CJ)3Q�5 �7]�`_�R�on��&�����#����^LP�P[aW��P܆� "���F�p�k�Q�`��FK܊�«�sl6Bb'' T�Z[!�puvj��P#�сF���%�������l&/�͖����� ���͵T�:�Mi���C���l;*F��=eC�s�7�	q���/�BJ�[C�L(��|>�(��p���9����Y�j�}�]��? ���vB����^��_}�����p ��+,X�t�F��,n�Mq7��ݜ�$t݌�Ø-���;��g,Ɠm�o$H�y~#4�H�?PR�/*�9���M��Q.�II�?��kT�-�=��J���Ǐ��ˆ�" ��B��]J�T�`�r<ż�U�WP��[��t!c�p�G.��:��[6+�,Ӷ6)����u�lZ�L9t������"\��0Q	kJD�g�2� M��+�u�#X����~��М(��&"\�Ӳr*�Fc��^hgh]�H�߃������VQH��+J��>�-cF��	^�-�c��}[
�PB��O}J���33�RA�!�=�����W~�:{�?�)m��f�.��Y,��u֨a��D\d :���9J2���)���~����Ll�6�D�`��5�+��!�M��wS�M���p1��;�3����(3B�s��)�-u���o�-�����1�S ��Hw�u��2���ݻ[6�� ����o��d�Yd�a2���A�4^�>Bi������^��W�l/\ @���0bSP�
�M�q�R�Xf�,]�D؎lZ�)��KA�[�4|ggWGT�<��W_��&	`)hjh,�O�87i@5��.^+��c����?y^�V�B��+_���i����Z�:��_xɕ��>��7@Ͼ��{��Ɵ��VбS�,f�xw��S�
D\;���D�et��`
�ֱb���h<G�k��2@��PON\T3©e�@�l��l��eͅ��u�2R7h�6�1)5+��7���Xx7���������kht���Lx^]�� �8�x-��l���M�KJf7
��:�H�-O�#4��'�؁Eh�`�h,`�><��`2��,'��0��Fc�"�-����7%AK���~��vim{���U���(���K/�ϞQʠѣ���M��L_���bmL���S/��*���\�@�K���t�bz���wz���e�e�I���
[�~�R����6�&t<-(1BX,1���g,� ��"��"���W\�Z ���̦pf|V�X$�T�h��㬹�1���֛���ECl2J�����#R��"ߑ���ɨ�
����V���?zJ(?��>Cw�y��\�r�sK~��'D�QG��bcx@Ƞ��i�\]�bvĝe��@LMN���j�~��[��fS> v*�eF�;Z�,+1Fgg�x��,ͯ~B��)|���H��� �q�e��"H �vP%�y�X>�@�,�`Rq���g$��|I�4?<��Mߏh�{[�o����oS�+O������>I��3|��X��w�N��{E���AC��PƢPМ�MfL��6�Jz^�P��r`A�9F�z�y�}fS��P�L�Kf�����M��/���h=�G�I��Cu����@i7M�v.14�#��׿�uY�x@�JryfZ�x��t
�{>~��AY� �D
�'@26^�%s]�d�b�=��%�����E�B��q�K���h8Tp �A��Ye*FN���>ѼР�^x�QI�Q)�'��ȸ�_�K�$oV� ������C��x�w��7ҧOi'� �aP�8H>� ��u}��/�W~�kTc<���y�~��41[�X�b��x���������SR"��%��[k��ݣ6Y�x�s��@*�Z�:�>�ܴ#�d>Б�C�Ń�'��H�$��7 �բŝ݋�?�݇�曮�A^����j�>�K�7��փ�U�H� ,C��~���i��s�3���xˍ��3::&�D�j��3	S��@�`�QxL4�)�$�hA|>�Η,],\�� �VD�!��1��6+�ா�JI����a�G�p9�*�l�H�����E��hU���^>���!�m���� �C�,Ϩ����?���I�ҿ�*��o�k�=��s�����NM����,R4Հ:��
1�]�՚�׉��Dr��I�I5�� W�v $D q;�`�}�2�O���X��PU�����=P���&�*��A����<��~��w�$�s֬́:n���� �i={j�����Ă{�O��OiͿ��;�]�~�$��Px��� ��^�Q����T3�B�o	��w�F\ s�^�6����L����[�L�PT^�}�C*F�6�a����%�瞳FJ���1)�4m�l~�=Ѳ8(2�S�]�@��$����%����0H�2z����g~B˖�����W����v��o��C��s/�w�K�X��Y֐��d �XJCI�����~�<�q�<G��N�tV��g�?��q��bY���h�<�J�@�%��ʖ%W�Q��0�5�����xL#��d�g1���y��	�O�G�\z9k�;'@��� ӏ)V�<�,�X,��O���+Ec�����顇�Ο�.�T&E �TAb���B����������0B	�|I�4j`�4E" �G@���i�jW�m;>��(�9l��N�V^h�x2)1C(RB�����RH�N^`�;�Rch�;?v���$�/�`��d�/_�n%|ƍ7�L|�W���on�������S2���n����̖�b�dn�1�$/�1�+�V�c���rϣ�kC�1�C��B��O+X�ua\g����ɞ#'U��יv�sf�h//�H��U$�@�H�YUi�Y����;d�prrVz���;N��v3{4�
��{[6�g��<v3�Z�o8� b���4c�we��⥔��g5�ᣏ��?"v����֛�K/�ӻ\KEx�g��":#�v"��ݩ|�2=�V6L(N-�P6���gdk���<2���6Z�t�R	���@�hh=o���<@۶���!���F1w(t�w-�����B��g�텃rk�<�oJ��<D�|�5z�G�R+�o�����>A� AO����|�Ƨ�8ݬr���d=���e���*��t�����k^��� ���S0��ǉ*ܻ��K�Wk��]%���C�#D������N�%�ڇ�����|��x��ϩ^�Y�#���b6E>U1��O'N�m��D70�B���wޥ�G��37)�'�nB6jlJ��ˬ�����[�#Qm�?��4%��{��Wh_��\�������C��R2iG3F������G�2K*�1������\:���&'��M����"X���eCAk�d<�^a���Yf��P&s����9�����<^~�Uz��'�K|����
��}�6\z���?��+T�Ts3�e���3���`"�-$<@�:y�
�;��QC@�qڬ��B��	�GDb�nNͻ��&�-�'��$�e�ԋ^k0X��e���袂# q���V��5b6�_�I�sz����q��^��ֻ��K��h��ߠc�Q�����B͔�Q��p? �b��?/9HG:!��#���_|)���
6}�3
���~����)thr��}�_����3D����a�c�B����F.L<������Lq0oP�Y�s�l�:I>���n�2�\�`X�<�������#�B�\'}����ٝ������o}�z(�1@U�-��s��7X����5tMGm�?Qƅ����{)���9�_^�R�XRw�!�gp)x�Q'����C���@��v��7��/Ȥ�Tf����h*=t�=��c�λ[���u�'���(5�_yUZ׻:r�b�R(��u$D�t4ZJ�B�"@�d8��H��G��t0�NG�d�!4��ڹ��瀍 ���@ٸ����T���Qq $�rB(^��� �c�R�����+�0��u�8����w� ���lƑ�A4��Ra�>~��|�u���'M$�����O~�6\|9��Gz�����tr�@]}�¤ɩac�y��*H{D$�*�vec�O7 +��M������+���^Ε^��*�*P�+poF�тߨV\�z��Z���	����]�h��zy��8L#c��4y�Gh��}�}/]v�G�^���r9�_��~�tx�)�aO*�*�L����.$����)�+ԿLm�AL�H*&��**
7��=;5vg��0x/>�Ρ�C@�����D��1�.{�C������e��HǻAH�wLŐ�
��d��M�����}�����>J��e�x5�ɟ�g:w������c����ǉ��:bv@|OƀMu>��TJ��O, 	(�'(6 ښqq�XҼ����`����؈g).���+��~Ih�DT
��-��I9	��*�t�Pc]��k2�Q���ʬOQ�Qe`?26K�S�`RN��A�׭f�t�4����k�clF121��	_*.5��(�_�P�T�QZ��?����5�ꍪ칲#���������Ih��C��%��e�O�e�P�CAB��	3�i�:ILh�V�>W�7�p��i��$?�Z
l����qߵs�$�����-7�&c�^{w=������LF�k�r�K��X������ 0숴��?l	'�
V��k}�H@�����:��i{�`	ǘ����A*�Zj�uZ���&�|si��:�d�_�rT]vd�R
hɲ�TgM���	b�kbw�Ta�<G�cǏH���k��}�}�_��W^�=���I.B�B�dP��� �7���X�o+��3ԏr�G�)d�)eԳ�x�&��8��M�vH̦97zO	���S*d�{tߠ����K.dsw�t��1����$�b����W虧"��-_E�������'s]�����η��E[������cA�b���.���*_�
,A�j�j�mZM��n�N���������Q~::�ԐN�H�+��b1>�����R�@��'zdO����x���bZ��_L��X����emƞb���5*��X99IçjtΊAb ���]�g�A:w�*��+����ϥ[�Y�i1�!!��悳`Yq�i#��0j�:/x	�}`�|~@�:Y�C�E`��[�,�UwbR�/�t6�Ӆ鶺v��`>{�z%���%L�В%�Q v�3R`��m�z���->@ř��R����}��+h٪�h{�O?����kt��5�B���S�-C2�I�"�Kܡ��v�Z�P���Q=1����w��u����\mj��>tjg� ��M{im-x�@��D��߁�H�@��h]�G��`�j�8!��z�jr�2�Z��z:��/��{`�q@�����S�3Oe8a�I0��������xW�֮^EKhl�*M�>���������=1oh���λB��'0��^`�)�=}]l�V�P�Vq��ӊmn����|��aJi4p�i(�7���4ojY~m�Q�>�\t��8�<��!�x�1��6�#�	�àiׯ�@��::������o~�Qz�'?�]�OR��=���Sy�ݜ�O�5�OIO�	]�|L%���r����F�4�3��bi�[���H�o�6ޠ8sl� 8�`�b����2 S/*�q��8��v\2&Z�|��8��4���\y�Ŵv��`	�ȥ�����
��ŗ��-[�go.�'�e�U`-��wov����j���3�齝�w�qZ�x-�.X%\U�����cP�!���������ݾMZ�+0�$�BS,�Tv,�<=�]�:,K(gy�q���v�x���P�*�51
�c �_�j�$�����$ݐ'O���M�+1<h8��ӟy��`-�t�8��O�ˏ=G＿���9�p!Iپe|ST��Mcĉ�g�y��Ii}l��rM��]C��l�w�#�H�8&�@N�i�3@r�̦0�r}�u|��-.���a3�m5�,���r���n�/cTh`ȧc�#��s?�����A��4�ul���i3��ƻTb��X�Έ���-ÛT)�gW����Ȁ%4I����l�ƞ�fڰ~5؅RD7�n�?~�A�^/ZD�֞+4���wn�139%�B�D��9^!P`Z�Y��B4ա���$L�0�T3�]{���dd�̘>��P"�9N�w�w�&ݣ��^#<��|�����hh�@���N�O7>I�����}���G��x'�Ѧ�׏u�lpT��1�:��؀j(��LI��m�pA���l��V�eM�z�V�yF���:��b���AVS͉>�
J7���5z�<����*��ӷ��u�~�n���i)Wk|�b�n@���ㅫ���\dcb�dV0��
k�����˚odz�&���6m�!�tW_y]�ћ�a����x���k�B��#Χ�\|���EC��b�q|6# �(�`��Ŀ=�́�u�SV�dZ��HG���[��jh�+����9Fp�!�(�Z��ֱy�������l�M���M[���쒉��� gz %�2 \ORZ	W=V	
{q�E�ڵ�"�?-d�4@���&���j40Y�
�ڡUc)�:k�/L�ި�l
#��M���Uh�e�d��2�����K�l�o"���+�c'�Le� X#�b@Ϙ��I>�Z��X���6��E ���_���J�i��5��_&c�ff���#����lv\���@�_r1�bp�I%%O�h��ol��t&p`�{�0h��!o��)�>@42���)�J>)�NJ+>4^��I�j-�Y	
_{�e
�Y���c5>1Eon�C���� q��3��9Jt/%��}�sT�1����P~ႂq���H�\#P�tlQ��<��}l�v�j�B��hᇡ�3�� ��
�K\a�%�*H��>�Gh��FR�3@O�-T�L��t�`�/��_/��1k�	6i ��	��P��Y��@���3��#�5%x�p�cp,�4Q(S.�E]�>	xb����=���s/n@���fՊ�t������/�PH\����f�hxd�=��7���Zq��Fr�ֳ2�%!I�����'�	�I�!9��=�&n�/?�i�l~��$����k0#(In��=d~=p֑
c���2�'�
B
V� �hT����.#[kb��,��(V���0�m����J�εШi*��F2��Eu/�,�)��K��E�B�jo� N��h�ň�Z� �<�HLWA,�ل�Z��%��������&M�!�Q��s�`Ap�����{��*�	X<�E3%-�Ma�4�\��!���mC��m;��S?yA��(�Y<�K�Y���%�[���>"'�d���xC�7�Q2|�oW=E��Iw6"
�@8�g�:p�(��O���s�g)ɂ�Qm�x7�/�j�J�'���Ћ((��!e������m�тƲ��,�2�5�$s�5��	�e��0U�V/�1��9�wX��{�M���+�8�#(c2Eݮ���M:Յ�)whU��ř�o KOLL\Lrth�b)�5��'���}!ocE~sa� w7�JUGpNx2�LbL�H6OB�L��t/oU�vY��&͜��K42y��Q�2	�@A���� =�����9T1=�$�H"�HyQ��P�R��(��)�� (�{����9�D�m:)�k�CF�ŜH�hPו�����VC��,�
"o.�b�V��;tf���lTc�"����z�RZ�(����z����sc����HWD�)�ы�+�1C�
�aC]��ɍ;j�bV)M+
���@x㮆(�g]�*�sI1�Y�@�]����$=��#!�@LR�� :��X��ޗ�B�d��M���e�M"M������:��&��� �[]������S?�3@>4˙�a(��>�H_(�R��y(MX#�6�@����mf-��i�{�Զ-�KQ��	V�i��c�E�,G�c��Vk(�O<J�L���Qzd�qq��6����@����
Q6��:T��U��:�0�A�Az]s"셶Erm.�����Fo��XF��X7�PV2(C$���O���H�'���2���Gk�*l�3r ��4�����6�q�9GA��%P������S0?��s����9�l��7���}���H��(ᨖm]/��9�����" ��Mm5�w4?7}���k��:0n�D?
���	Z�`ч���.X1?P��]d�t�j�9���� l�l� &B������.r�~T5�FR�ࠍ̋���C�9�<@ng/\�N6�U)Q��dxg[��\]VA0��V��
�C���7:�ZB]�-1����O�u���Q{T`-Zkpt�؏R'4�Vտh��=Z+=$m�4CS�E!�=-�)!�OP���h��8go��p'�;|zS�y1\�/�g�$3�MM��m��\>��1�VO�U�ZAakV��Hf����zU�9�˅		�"a�bosQ_'�O�RP��I~>���N!m�3�p�sk��-K'C�p:Q7��wC�/�j�B1Q�����x��R�PȬi�l�>ڴh��6�b��vϭ6��XH��c��j�-�{����k9��y��]���O���zz�J!,`C6�T4F��so"�@���dOm{Sk�F�*ڄ*l9q�9<���Uv���)�Y~�'��<-b���W�W��I��>�p�'?a�D��?!4 ��#ω�t���&�تn�z]csB]'*r4p��p��1i�$:F��/bq�������&�����4U
��{¶���|n8/�M
d�Qўo��Q��QK!�c;�b��4�F�����LIa�<�@���t���.�s��pN�;+\1c"B��$:�������_+Rif��)�z�Y�c������<�^�\�><���t��1��i�f-��t�MNI�H��8B	��hژ��&��rԒ��i��d¦�R�����y!��r���9�v��)�w�N�- ^�,�9s�N֦�;#�!�;x����KZ�����迖\�fUX\��5�i-�T�8fꡬ�ͪi qިDuX{u�y%�FeZ�Y�{��O+;st�G��Sc���KoR��X��4�ڂoBW�}&�`�sM��:W�6�#��f�.~x�� t\c�5(ڲ��i_�
nSE9Z�+	���m�rG��i!�)i��8�s�&�E=�&���Y�3�9��5���/�?�`���͟�@\èvj�R{
�
�0������i,��gj�����0"�h�n65�T���~��ˣ�Q_h$SID�{��?B���e������s�^����ݒ
�\�ݫ&J6��1�m����Kh�_��>#������m>Zq���[ׯ���7Z��������<<s�}.hoj�0�iF�U}�t�K�zZ��:����`�%~�/ ��m��N�<!k�{��k��asK��՗�ِ����$���.�V��#�S��ɟ�&V�6�iO���G��:���*&6�q���^���s���>J9���3�3#/Rs�ڵd��ܖ�W	���RQ����h�Ē����y��B�{�XX�MPs�Wk!��w2�l��皾���4����z=�+�OǊ'�7�V@�N3���`����p�Z����q��	X	U��.��FM��W]'��|Gtbx�܌���ӆ�����)��	Z�}^b:dx<�D	O�@�wgLlTK�@u�9��x��S�����m��Ń��B�M�Õ,뭪BQЏu5ެ�~<b溭p5���$|�f�[�371g_��{�W�^A���B�2�ªV/K�ᶜ��mo��ʌ�!�J%)/I��Ck6\B�׬���S���LwyD�ӛo�+e� ͨ���l.�W�p�K�#%jC��6�k<H��׿;f#�S��J�L����u��v�x�=4�������D�Ɔ�Uq[LU�M*z?&�᚜kH2ĉ5��Gp3���Z����{c�$��D/+���
��4SJ��h-�o��ӛ�d����-ƴ�`E6�)� s��B�غ����߁&T=�.��>�?:B;�����q!	H�����MO>�S��8._I�l������aҰH����Z�F��\[KW��h�+��P=KI��?����ɵ�.�hИ��̀��������������.\)K�k�P�N�h�y[p`\S�e)��vDV��I�ޭ\�Y7�����ؙ1��2-�b��y�*\�V[Vw�G��8?l
n�Y�_�3�[��'?��R�D�>�Sںs�w�Z!��w��ڳ����z����b�Ɏ$vØpl6X%�u��F���X���U�sX�s#\��w�Ѓ�/n~��6�2�KB����hdH���j&���x��$)v�Q\h7Z>�k�p[-a�و���s��N���� �Ms+0�Vo;d�0}�^�O��ɖ�g��/[DB�H��h��������Ys��
U��E��u1������x2���A��E�Α�,x�,@j����+�RT�T��t� fC-����uv�<jb�V�z��=X.0�:������-I��B3k�/~Ska,r&%�/�����c U3Y�fC�uFĬ�9g�`��h��&��*&��C6��b1�D��XC;��.f|~8&�����x�V==xOWs��5����8�ltR$|���6W�E�9�%d�9��N���4�%���'�)X+���S�[��)�$��i���{I��J�$��'24fBpZ�Æ.�uV<�R�Dh�ɷ�L4H#j,i���#���JU)}o�U'�4;Es,ضo]�֘�{��#��u�>���-��QO+ҙ]��V��\o\#�q�c
˃��i�C9�h$N/X�t�l���E%(P$=���3?Z�-g�Y���0���S3i��w�J�g6��fLdfb	�����:裺R��д�i��+0���.iC�Y(ႆ��R��j�@�
��j�b��'�^��C'4T"fds�"?�aS�����`XA*�$;�ıB6�@�h)k���(�g,�/���`5��@jV��,.P�Ύ����&�覻�3T�d*XZ�~~�tU�F�vz��w�(���@]���Fm;��RB�5�(���k����>\g�?6�26���k�vL�@p�Q�Rd,|X�*5�&��8E3I�V���$��6&D�TS' �0�-�!���S	�g��#����s��\.O~�L����)!�ŀ�reJ�0b�u5.�Sꮤ� �Z���\&���D3�i��9��Ñ��IÈZ"ֶ�<���5��E=}VPb-pCㄾxrв(_��8C-� ��W��5!��~L=����h2Τk�30��d�'rDm�R�#�
�j�zz��/�qt	�b5�x6,w
��ހ�Np�4U뉳3Ws����p����ba]����%C���e�c�}]����,XU�e��>�8���WOOLR^:�C���{���F��2�eS4;r\��vK�F�� /^�l�ě���'P-���>ũ	�9+|�y���嚪A�����DJ�M��X�ԯ Qp���V�4�9r��9��M�l� 0�[�bc����c�!k(�� �-j0��>S��FǙg�ک"k�� �7xm�֦���`��67Gx�z>��{O'�ss?�>75=&�Y=�G�)O�����'G�������/����'��-�Ks�4SP��O��?g�39z���7z\����0u���s�Mt�5WS��bZ�l1�0&z����M���C'���gV��b�l�X�Ăg8��ϯ]��n���󶛵��Ҡ'�x��y�9�(�ױ��h1B�qrֳ��V\e�墷[z�P��F�%r�`(<U��tZY^��Gy5)�ĵB嶘�|��X�m���:�	GN[���*X��3>�vv�t��0��y��¬C����ZHI[af�:�)���:�̥x�ج&b4[)P��k��*��x��)vx��R�r,t���_�;��Q71��q�L���n������7���c3�� ƀ*��5v0\ntB���c�g��`�V�����͎��O_~�f�c�L�y�i�dR�|�o�g��ߋ~jI�+��umD��:���`B��)pUqd��q��M\|�\W�`-��N����۠}�?�`ѡC�D�%M���F�O���t��w�t�B������& �r��6	��P�qgQ�56z��ѕ�_D�=��!�W����brk�i��u��a/�V�|>CW]v�u��Ԩ���������?�t�H�V���}�W��s��o|����):15+�6��Xg�7[lPcz�v�)���^>v�~���izj���?����~򋟧���B�d'_C�pC4�AJ`,�M)[E���4���4_�"��{�Z�⹮��m �!��k:Ѿ���sea>یh���!�z3�M8�܅g�]�kN�8�{]e�s�����G\�K��0�m[ާ[n��M�-�����Zf�Wa��}Ǉt�%�	/���/�d=��Y�ds������}���	������c�8]�����^��FEkIZ�X�;K�C���u
�K�����m�K��B�'gg(�ꖆ�f^�9Ip��,-<'
O�R�ì���B~v��]R_ґ�M�92�
=2O�����h�w�kj�ӂ8���n�)����������d�&�%ο��a��@�Cg��a��_��k��B%��S��u*���S'Ghld�ְ�������^��+��c4ujZ�xeE� �ӆױ���[�b��c3���RU�_=>B���s��� �,yZ�<�̔��,ߑe��K�z ��5���߇�:�7{�i��-]8�L�6�(R�l�y��*�#+(u���w�n[�C��Z��v^A�b���06|cr!p1O�"蔒�3@bn�8����3��+��F�?Q����a�iZ�+���5sź�$Dg�j ��e#Lz,haM<&;�<�l���g%]|�E���Mt�eW˼�����ĽɔP7��V���w��)�f�C�3�S��Q-�*��J�H�4�ש��^�2�$}���Ӡbէ��QZs�
���OP��ГO=-����׬,�8��tט'q-�j���ޡ�ٌ�B�r�U�����k�����ؼ�P0y����f�W��4b��u(� ����9��s�)Wy�����h�v�D-�AK��
Ck��"�;�s-,<��([_��;,�cP�����R9���p���[t�mw	����_�k��J��ko�A��N*UX�ju! ��
b�$�0�/���_�W�$����<3��.N�t'eso<An##%G�F��k��E����7	e��қ�i�ֈ=�Wi�HPl&By�5� RaK���\�^x)���SCն�(�����#U�a��j#�i���X!2�~��4\mn��gE��9�i�Ӏ𹏅��\�9[��Wџ��oY|�L�øaNVCxLQ�f�j\�K�ןG��Y:6|���2��#D�Ha�G��B����r):��\�ԐH9�]ݒ�9~�����޿�����(Ş'�w��=��OC���#G�)#]��{���4�q�{~�A�m��v���キ�f�u3*�ɵ��,���JƠ�ֳ�o
hL��^�hz�c>xg�q.Xl�j���Z=2K�t�c�xVk����ل
�O��d �dNrqU/c,l�jM��Tm��h͚Ut睷J���g����]<0�1p�=��G[?�M�_{�x����OQ��wh�*�Ӵr�b:w�j�^!��s�2�n>�I���X2��Y�Xa���q��������ߗ����`���y�P:�fp�hYU�4�4j�M�u]V0袲�9s������M03��4�'�q�dUG�Yd�_ۼӱ ���D�m���Zk"���)�$�n�B�`g�ӝ��G tDȹ!�T*ϰ�I�u�8B�332�TH�ٻ��߰����~ؾs���t�`Zh�9.�7�~�.��J��o����6M��5K������&n���,����|!���kJ�7�-��;Bg�ۓ�?��ߧk����~N����Re�T:�\��/'�_x�%^4���z��M�|/r!h6�%�1�Ӳfa��e��]Ȭ�g+�[��r͆	���7,t�����?�5�g��Z��q�@�}�f׸��c3Vcͣ�Jt ���D?e#}��O��)Vh�P�͑[���)k�*l �;����>{����˯����RL+pbV�"��wh���B���&x�lJg����}�.X���3�t�5W��\�涃≜ԙ���}�^|w�Bl��svҒv8�B���K{��i�V�+`^��ȕ�?����?p�ɤv�&G� լ��c>�R:�6{�J�1��`Q8O ZU����羧�;Z�7h��J���>Ֆ�2ǅ�!�bO��Fr)�22*�B������?��&&��:d��]�@��r�ƾ��th�A����К�k)��h߂D������[�Q"7@�����N���D��1X'o�r�>��������N�	V�N��@����N���Ƃx���]�V�aٶ*�5%�g�o��y���>�_5�S�b oݶ7-d
zk�tt]�x&����W�6#�����)��4S�-�`ӕ�wH��'�R*��r�H����ѷ��;�=�<���X���?�*`�<�?߽X���������9��MH��ė���{[鵷�f�hP�A�7���A���;虗^��Z�T��5��VXk��c4S���}�Q���X�e.���	��Y��ML)��"2ڪy�6%s&�X��F�O�E�m��)d*�9:f�C-�i�8+t�a'S6�h$�,��3�B�̧J��+�0� ����`�ߔ!=�F�-��]c�C�mY	�w\�߶PsL^�����lZtI�
�B��R��iU�r�dC�S.e�i��ץK6N����<��Ta�����)%�`E6� �-Uz�ӯ<�YZ�v-���HϾ�s��֡≸K]=2� ���K�5UX�Bf;�V��+�G��ǂ���J�#��}
Ȗ�$b����jy�,m�˵e ��4�Y1�h�	�xU�!ē��Z�̦3���,�0��B<Q5����^�i�����B��8�hv��(�M� �=�u@62�\%~����hF˘M=,�S�v�h��&h}��oA �x)�AJ��x��{��� �*C���ע���s���|��l%�I�n*&f�%y3��C2ɢR��3/l�%+Υ�����>�ҫߠR�Dq^#tl7�x:�Ԓ+א .B�\�/�`�V�C����aK�A!d,pl���	����|�*$M�U���qYoOL��c�ʳ� 0pj�q)Rb	��WA����ar�@@���8B��V�x�~fS�S�l��KM4�lh�R�H�j�CvaT�i�dǉx�����t_����Jhs A��&l%v��8�ś+�Ԫ�Z�I�$Ϧ$�YX�)P��xQ퐁�P[�u��Ed���ǿa��.��@�|G7�����?�?��7yS?�y=�r�c^BJ|3٤��&���C�w8qdn5`�j����>T�Z��j!k�5���A����f;��oH 9�L��j�D��6p�"9�M�Ϊ^m+4Q"�NX(�x�/f�Q�!���C}6�Վmdp�u{�@�>�Q�+�|O�B��Q�@��Y� ���ʅ7UF�A5��T&#5Ldl���1}�Xװ�o#Za�\�(�6�Gj�K�^�(�c�^�_II���|�I�2��Ԍ�3`ҫ$�;�3d\.�<�R��#�U1G&��q�{��в��;<װ����9J�P�Y�#q&\��
��N�H�M�@�L�/�ɣƶΐ@�L��~H����0,ȧ��#N��uvW2V��R';5����YrMձ��!/���}��^&�dh~���<�K�k8����6����$��ӌ��4��>K2Q*�?�w�*jÑ�l��dc��8
z�ۢ��!vj��[�IF�8M��Mϵ���	e#��lrrf*����9�L`l���K�B��9(��C��R��v��H/b`ۯHcEdU��A'����m���35	N�m���ݼ�P&�0�K����Y"�1�@�l�'��5�b�^PڣN>(Hke��J];�j���?�ae��'�a��ę�a���b3Y|G3�iV�H�V1�/$��1|��_.3�@p�D�JIf�)�m\N.Ʊ��s^P/��,��@
�j����E@�3^م��S�,9ԍ��F+T*d�Vf��<��EF���V{u����D!��L[}(�<!Pr?�]�I�,�"C�`��C0p �Zy�#ѓ�4y8
[ۻs��	B��n���R���s�����*\�T�h�܆�]<�&1G�C�OY>l���q��R��cy��:)��&P�g�=��]J��Ar��0��pc�����$�g�����EB��&�ǟ�F� �F=7��um�ʲ�/�[̦#!����t�`@���%��Р�
4hU����Ϩ�߶9�ބ�Iq�XVB#R�L�0�Ykޛ��v5���I�뢒�m�B	I��<���	tؤ[�R�q#(�-�
�4���ze�	l:F���6��ֹ^30��C�p�P�C����@k����t��c������:M����QJ��|�"��[E�])�ݩ�	�����]�%�֙x�Kg�$�`9/ҏ��h�%��bU�T��/�0���k�'����5oԊ�fo�K.��.�������2�����ct��0��}�������k�|��I��|:�a�o���:���  5�IDAT�k�e�<N��\�1&�H&2':!p���5	��e�	M��1��k�q&�VB���;�{A��B=L����J�����Zi65��(�Fk��mƑ�w��Hd��>�
ikWh����/J��ʳV���R�4A��l*�t�W�}��M_r�̼��YFo�`�]^�C����?���cz�w��g9��C�{�9D� `��\1X���j,!1��UJ�gPg��ڕOSw6Cc#'��t�%�ݷ�B=]2�avjR�.�@�Xᓻz�-]<H��/������Ghrf��_�Un^d�U����W�q�CN��W͇�������-�VO��73��u��B�θu�<�Y�*���I0)&�v�$�	BS�ь�|R4[`}���TJ�ݖX�c;��a4��Kٟơ�y��Qu�&�u�e��ϲPud��(OҩchŢ~����7]'�15v�
�޷";XS#$��7��O�{]q�%��3/Ѓ��*��1J�%x��T���݌�1�g,�s��,�W��6�#�[+��P x�u��5W]B��;�Z���R�p���bZ�4`:���\ͥ���E�x��"�Q�^�.W�6�̢��z���'�&Q�6@iDfq%L!J�+�����F��aKC�@�O��:�Ơ��1� ߋi�6��8[�/�I�@�{�(;��7��VrZ�i��j�U�k�ϣZ+�1�Ѓj(S����hҖ'�:�"��@����-�h��љ��n�h��!Z:�M��o}�.�xՋ�4Ç_���>keG�.�Pf�
����}���~�kP'c�o?�(�=r���:���(��V�Ĉ�$K�B[��<���=_İ8�
�b��u�`���\��ןGW_~t��k(���a #:se�|�(h�g�����^����[���7�F�2k�4�ϘN(�#Nx7�j	j�b[ m �@�t�	����5�n6W����i��R&Q|^@�JY�IO*s��w.1:>�?"�Ё�!GCit�0��`�)������r�B�a��'߼��<��8TL;�a��$�$#i0&^c�zM*>C��f����z�b��'>F�[I�G���%0
�4�Qu� q�o�Y��da�Q��C_��=r���Ϗ0�9B��&�%e;�T�<�+���1G��ǆ��E�AШPw>+C�מ�Tkh<@�A��c�Mc�,GP���[ɂ���th�|:qd?m�u���J�bґ�ש�fz��`"m�P�x6�������9lr]rh��&�9Z������I�n`i��5�^�VԴٮ_��ɾv<KT���0i��Åߗe捲7��	[ Y��|�2(���a��H�#�p�̰
~�������)ȥ�T�'ׯ�m7^K7\{%%����Zw��e�E(]�[��.��#?u�mt��1z���� ��Ĩ�Zc�u�o }rf��o�u���d3	��$���������ES�X���&pb�hCk#������j�N����5���Kh��8���/�%��:�v#m��M�û뵊�,���З�Hb7�E��p�r��+����G�Ml8�!�x����� 8�@ӆ�aD�j����t�4d�J:�P@�b�1�P�Z�&	���QD���q�W�1������޸#��EGZ
��Pz�F]&5錄I�*Aٔ#����h=�����Y�<�|�1��S��iF���AmPA���T%�^C�v_�ґ��i��s�6�2/�b#8y�������g��g�X]BP<G��$�٣�g��%�e8v�0&�ñ��U�iO�I���Ǥ�AǗ��]�X2H+W.��#{x���S2�8��:#&4 �1t��LROf���{:|	9���A�0���S�j�GT�i�2B^�t:.Q���tT!T�D�������13��)m��" 
�>dٔs
��&�S@ z��K2����$Y��Ų�%L+�?���H�U�*40���'f�H�brP�(ܠ|�(0�#P��/ѕ�������C���l��+fLK�N�@�����g�.u��ʣ(a�K/:�n��*�y�u��*U��vW(D�r=g,|�-��!'�O{}=,����IV�劘.9G��0$�D�7�D�e�;g�,�|Jװ����>��w
qr�(s�(���au���d�����)�U
�_r�T/�x1�,����$3�ꗪU�/O`�㞉��)��׸hE�I�HQ��\ma�Ch�����4_Ogg�Ҭ�fI\
�)�3z�;idb��$�'� #0���V�X-���,)�X/JS���C�;�q��o������CR\&�ńg� ��Zxb�~�9��B!�=!I�ȁIɬHm�RGZTH�`vk�\sB�M�Y�5kVP������`�eBY�e�{fS�����d�Ɓ���g��<����� ����+M�[��~���|�����#3|3%���Ӊ+�Ib�����
���,�� �O(W2,2p��$L~^B�"�<���d���ŋ:y� -[���;�4[�H����2$s%S�h�L`�L`�����5:9"]�ld�O�=�k��q�J�Hu�őb7���8d���ϫaZ+���)�f�ba�ǫ'�������3�|
��2�:%��pH<	�_�b��@�N�E ��y��*^x�1)�7��<_��M�4���С��5hӠ\��CaB�2�0�9K������F�I�͠vӌ�j2�����H�x�5�v�2�)+�`h��ʤ�S� #���ϔ��*&��ڶ��w#����3,P��a�ki���ɉ-죎������O��x���}�92"�y(��Iu��d����i���t�9�dP8Xc��=@GO��_bӔ�ɩ�g��MVxA|��S.�fYS��e����z��!Z�t��c�!���_�Yh?��iI6''�5)M��k�ko���[�������]���C?N�������B�. ړ n�)O�80؛n��,;]%�>8�	�·�E�U�qUCJk*��,-y�sb�x���t�����˳�vj����!c����L!�b?�����Xx �|�=�YZ��)Eucc���U9q3/�!&YH���L��τ2)Z�OP+���MG��b�B#�Z0�a�}Oƕ� �a/-��e}�R�șhQ� ^�j�q��id�"��V2��b�*u`]��l2fƎ��(�`�5M����d���������Wߣ����� xeV��OT���4����1���~���z�MD�:Z���75;z�v<�� ,��zMbPY~ry.�K�8N��m8o-]z� o {\c�����=_��n������6���.~����}`:j��5l;>�1F�a��H��.��5?0�PL�T�k��p?4$ Af,�d"M4a��bh>�\4����ET������txF�����bCj�E@�Um~]&�g.X+C�Q ����BY��b�x^�?��"�S3Xō�h£�=6&8!f*!�#�&�'����º���":�{���
5Z�l?7K�V.�����i����Ok=�I,,�.,6]��8u�^��3���H���c��;D�l8��{y� ּpɸk*6]��#�T���^6q	�Ѱ)�b5;1L�ޛa��fS�A˗�(�Fc!�y1����Y��G(��!�������$�?˛���ї>�E�ؽ���\C[v��S'�kp�T#�(U0�}������/�R�&'�i�P�ZRoړ4T��R���%a�)!p���*8ChQ�295�V��8��bV��NP;K�]�ر$[��8�L�zww���O���QqQ�W2�tN�(f#˨S��'�,u$-��i*1P�e��)R�Kb@Џ5%�>�ʱW�S%�;�W��8��R��r��V1^�3�}�7{u��"T8���O3,�1xAlZ�G�l���"ԑ��#��-[���%K�q�?|����&h@�?�a�,8��v=�&����<k���=t����`�������ALJ07����׎Ӳ%}��5�у{��j�9�ݰN����4<2F+�]J�]|>��i��Ka(Dr��	g~M�/._7X��Y��w��:�bM991F%^�T��.�W�'���奲��^���3�7ĥa�@�<9Ja%�	� '�֨{��v� )����T9b��!4x����8�޵��Y��O�$����?`��������I�����f:�XmС�'� n�\^�zE�����WM��s��R,0f���W,q�����N��=�}��}Z~k�Dw��lRf� L�J2I©p�9+��M���	���a�]���yz����g��}{v���s���?F�w�-��,������n�Z��M���T)�i��!���kyNһ�oea�fݖc-��S#��xd�x�rlV+�3�g�޺tު�2f;v�k��x���a�z����|].��6|d=��[|9Jgsb����V�T��|T�3��M���N���1�B̞%�8
( �j���?�ֆ%$����:�|��R|�����fK�(���"�%�b��g,7�,�TS��3�.�S^s�t�"u�d8��rN�+�=�&<�e����qZ�O;w�0e@�%�M��.hHes3��A�#u)�M"pY��ﲐ�VI���bqX�O�4��i���S�I��	��!Ց�MӚ���8�4q�x�'��cAYGs��0�4�}ϭ�t�Q:Ƈ��0{���dc@�r�v(����Eڳk']s���=uJ����u�f)��b;h�Q<x�H�3 �%�����c�O�	��_����IvZ�l�C9�Z���P�� �#a���l�J��=v|�^y�u�����t������9u�N��@���h<�<6����#�������{��~�}��f�G���6�^�>���*F�B[Z`R(Rx�DA��_ڠ�'O�}@w�vK�'��8p8��F,`�eȅ��g��ɧ`�ì�={�I��N�|)���p}�#�&��1Ʃ1�j`�/p__/�x㍴|�R�`A�[s������y�RbR=���/�R6�kl�=����iժUt��Q:uj�M2z�������ჼQ�5i,ߓ�8���S/���I��CZw��b�
�Ŕ�5:p��~}EO��J�V�	>��uhd�k��B��a�b��FJ�<���i�p0���Θ�ZZ��@2���J Zm�5�-[�������jZ�Xt��4�]��㣌,T|\Ye�*�ꋼ�1����C�G��@�î���Q� G��	��NUc��1���]fj91.��˨d)G�j�X�ڜ�[wP&���.��-�KE���A�q�)�ǄxD��	&�i��^�ݴ��ly�O�,�sK���!yka.is+TD1����a���2c��E��m��.m�ʋ�?H��^��-�n?N��J��h
�|�x6!��Kzs�?��z�D�����}�hlr�V����X 0�魷�ж=�X���v��$�{�K�w�KS��]y���������ْO��`��sqBX�:�d�
^��2ɚ`��A����hr|�S��o�B�7��Pa�n������&]3Y^wh�*��i��o�Ӆ
9Y�5 c�S��s/I	�(zS�<���)	[`�{,-Xc�r����b�e?J�>�z���tr�̎��.�,�^��
 Y d$ܳRo�,��p��.����ebIb8�V�ǟ|����G��x=�[�F"��J�� �` !ʯO��d��?9<Fﾷ�6��6��N�0�_ɥ5��0.$���
H�4�]e������I���~���;���O/�-ZNÓ:r�1�D�c2��pj��˦|1��݌ubl>f��^��r�w���;�0 �_��X�*2#.�$_���|�Yʲ)@����؉�6|�B�����KK#��of'
&�t:h�/ߡ��\A����+�}��H� &�n��iΡw�m�`�$�s)�F�'�`^��PRUq�g~�a@�2�x0��u��I��[輵�H�S���ڠ��	u,a�M��>޳u�A*7b����#qi����
Z�H��L��Z�������Y��E6'v�]���-�w�	9L�[K_t�Z��Ҽ�)�)���c���~:|l���Wq��	��P�EUb�|��2��p�C2�K��G�Jf�28<��˧w�b�e:�*Zɸ
�(Ϧ/�8�U����9��M/��v�RG�ϛ`�!��,_CY0R�qג��i`�_Z��g�}�:tl�1E�]�>�Ê���BI�I��\-�i�]zx��W������f�}���Q��#����-��ldB�+�]��CM�)��Mt>k�O~�n:�ܕ�r�� �/�������hbl��� �&�$��fԲA{�d!.��L��ū|Y�MM��ڦh������Uln���]J����lMPE����{� k��I��V I�.��^f��"웄�<Ӵ�Q6�����ڦ��4sƤ6���&��u|�F�V-c5C�l�!q�"�|�I�)v$e`���,�O�XMô�B�g�Z���ၔT�/�����y�h�,������)ӑ��)��ٚx���0`.�����Q�
���� ��E |6����+����������K¨�N�*-
iQ�?Z�W�
j]�
���V[�u��ED�P&��Ƞ�E�C�%/o����>�E1�k[x.�Zw%y������nJ�d3��n����s�!/��2�b�j�>���ԎAv�Ў\e� 4�g�#K����9ĺ#�(6ᾃ�I��P!iB15�Lĩ(51���3tZ��"����%S��L**w�o���^i���Ⱥ�[�;$j�tҡs/����$��#���w��j,�s��(@4��d�m���)x��T�cC�"4G����g1?����VHc<C4GŠ]�L>l2� �DoP��d�l��(ec(caPLRU�m1�>K6��Ҧ.��@c�	ˇ
���R?i���:���RҒ�HZu��AJa�ur�ĉ\�á纴��8`�ژ��<XP"T]M�:V؁�����X<"�E%إp��!E�w��0aJm�[C��ih�!�̑*P�kו�����+a7S&�(�R�W�s����!�,���ʋ�H��0��6�)�M��fٴ0c@ �A{ԷX�]a7�����2c�W�S��5A��]	�+&I��I0� /.��G��A�4��9�9��4����ąp:̡A[IF����Fʂ7�"����:���Ͻ�*c�`2^d<��G�l��gi�@ 6�o�m�
p�j�X����z���j�㺋��q��60K�]�1E��)*��	�X� �M�
��:����n� T+�".�yՈ� HǬ�̄�{����X�!f�Y.��
�,����@!\�N�H*������AN�D>�\@�����#�����P�hZ�2��D��Ds�� �,d��������[���8܉3ݢlM����
O#Q`���Mǁ!����IA�o$m�LZar^b���V�n��:Ds��?�
��)�f!q�Ͱ��ƟX���B��˧��0Q�by�Ȳr� $�̺�}��$lƪv�E�"k �M�a�f1)�2��#o�~�5�[��(ʾ�p;��x��R���2��L�d,2�� +�P�x�:�u8���Ĕ�V`�t��*��v�P�M�!��g�ƹ��AY�5׹�IK����3�3����I���y@�b����$n��<0�!;L�_�C��0/Yf�XI=�)��c1����P"��::*;�sı��c�%(��-fx�, kcy�/��	�e� �qrgX�E~�@��1	��t�k�u��ũ,g���6]	�҈%���Sq����-E�9���@���(�Ťa~�J\۪P����͌w	w��)C[⢔M�U�AL�b��0媋���$��gX[蜧��c�UT�:�� wm��J�eYa�d2+��� ����Ǳ�8VNQX��7�A�������b�����Q:l����F�e��j =_�U=c����Z*�Xl�a�Y�eP�6AĨ��,�,��CǄ:'�֓���@��v��z���suL	�s?Q��)�%��S�"'u���T��c���Fl�\�9ȱ2�Pp�&�+"�YO1������B�M�9n�2/"a�9a�9J[WZ�,o�zca��n���j���TR$�k4��i�q�t�ܳ9ʹ�|�@+�!6�J�]T'+A�h���הk-Hp���Ӊ�.'�졁��5�wK�2�G���ZB���8Tel/�[֌�ܴ�ց��̆O���D��0�4a]��p:�A�x�-$Rf6����#* 6JVf�S[A�!T;�0+q�X��صƼ]�a�k�4À�D�&��&BV`�����e٢+Q١���C`ɻ��0;��B�se�؟sDŻC>�����.��5J�zt1�8(�U�L݋N�Yp��M��\��d�8,8f5%�v7��L��X>�x ���(R*c���>��A�qEPZ���E���0\���<��ʳ&(vn��5�h���0>^`c�$��g�(PDQ6�'.N��V���\�pgD�3Mf���C<x��H����
,j�&h A�]�I�U�NVtLǶx�B(��D:��gT̝���\�)�4o$epb�����2�4{~2x!vV�І��@�"<PaL̰j yd�I`C�/�5�R��á��)VK��
��ayR�L�����Щ��@(�N,�����$�2�\P����T���A�v|xy �e&:���u�B%b�24�}��������7ޕ�c$�c
��[��x^�\..�GR��s�~��cQpf���d��p��'�ݘ2̨A�\�|��t{x�m[prnI"K��6���A�r�5���y�4�e"#��#l9�;�-���)�J�x��]�i2V��P@��R�}�6�L�Z����/K���-�i��)jC&����Π���m��Qjpnu�?��#x�4�Nw�P�Ia�DiP5-`��R�LG	�T��q��Z�`ٖI��'#�2�f�\б�����O�Bp�
,�M�$�	�piIj�?��h��e8X0��$����Bz*�-$�XU}g�Z�[�<vq�p�M�^��
�<�+�n��#|��Ǥɦ��`�	��`�l�M����:� G�$�%&�m
'���d��&=��a)uZTi2dH�R�{�����	������dHsJ�*i_}��m����%�ׇx��4�u)(H����$�I+WVD�S5g���ܾk�ƨ ����|C�s��������o�)J�H�L<�=��aYw�
���W��@0<td�x�Y/��M"�sZ�pa�7V-�7o>l��UW]1	^>nƂ��o�<&֔��c�vkF�q�l/�3lX�����R�ɲ���1�r��d���?<m��IpM��ۯ�QR�$�(�̰�D��l2��H5�/�����[�/������<1#�8��f�����q��Ç��^��Mh�l">P+���IQ�3��/��ڋ� ��z1gk!/�p����l��O����*g�O�����?�[�����F6[��+�&�$�/"yFy�XAY���E���$2�@Աº�⤋T&Y\]]�`��f���Jy}�[��P�
|�^�:�5��[���%qG����,��\H'�N���'���c-�4��x�7EEEؽ6
*:d�Z���a���t�kY^��Jy�X>E�8A�ܠ��ay�x�L�5-ñ�"7��IJ�b1�o8��<IO��q��1,/d-�4�<��g,0�4�����(U����2,�œ)� ��C<H,��l>�:3�aq3�L�du����v N4�=c�Ab�0����4M�$�0���\w҂E�Ѩ'����)������Ҥ���������qt�g���e!t�)+>�ݼiڞ����bY����i��yb,�,�Up���y3��9	&z�ЂF�򞱊���t��q�i{���`�w�G8���$mb|�#K�Ɏ�x����ph�qZ��䌜h�{��ի����np��izR�ǅYGl�ֻ,˞���T0װ3����ӹ8��q4�e�-
&��n<�����p�[n��FTxQ�,-O@\a� 0�u�cG�PK,ǛWh�����϶h{R�'�򞱐TUJ'9I��B��-�u��l��%l��C�u(Om�ޜC-�v����z��ׂ����@�����O�Xʈy7l���%���xZ�.(�MP��!�r8�F$�$��k�X��İ�R7�'��[6 e༬eq^m,fx��^BX�'hJ$o�$���@UҶ�?n8!�K�F6vI1���%l��놋}8ED�zb,�r�hSΰAzz�4�`�\��,Ii'�X'��@0�`�C˦tO�DC�����(��|4�Qja�ԫ@�P��2���tCJ�,�g��`,5N
��M�X��V�6�c��)���W�
�_��KaQ�e�tVa�;_�C=Q��`,9�ƆH����!qR@�΀6@%�Ib%	��(����0-dg�`�p^�'|ى��c	�da�5�'�7�e�65�2�!��������c�{szYÒ,Kpiahf�%�����IN�%3Ð�1A<���Ct�NjhBʛ*D�a"�Whgy�?eMQӈ����g�zpL򎹾�ED�۰$�7dۓ�l�fPWm��lb�P,x2��	| i0���͖"(*IYI�㪬7uk�g�q*��ߦ��
����.�h�
$������_��_v,��T�S�1���9��>U���]�.��VϹ�:;v�����!d�YUU�ڽ{��(���Eʃ�v�b5E;���N���K~������k�Z��"2�ݵwj���Z��$��Ҡh���ۗ>���9�Oc�Ѧj�S��p��͓�kMW�����a#�n����Z���;|�t�E��ܾ}{�����ɓ'�Ouuu����`�.]�駟��A��.++������_����«K������}s�M�o
��5��z.[yϯ^z����Qš'#�-c=��O�9�gU��ǚ갑*<�����^Ŧ�`նX���J�0i��wk�'��m��C��a��z�Y���6�6�2����ܗ����5���{�uۏ��3�<s�m��v��M�.�JI�z
�߿˸"�7o�}�֭gO�:��	&�o��}��l���߾Ohl"�E�t��Ui]qb�������7����o.��C�$��e�=�C�7��)�ٯ+��:MY'[��8S"dG}�!��ʶ��=��g%�k�W�[p�^�5��D"�D��-$b�R���*��7�ն<��r��޽?G5��COY�v��BnVM<�E��p�~
�P׬Y3޷����q�"nX;)�n�}Q�"T��;��)Hz6����D���7�^�:^˝�$��d�[����C�I��'�1i���>we�����C�~<v�����/��C-�[����^��cG���f��]���,�?	J�<�{S]v��n��5%��mߞ_-^�j�T$��^�~��7�k;r��gM~}��A�q0�u�]������uȐ!�˗//Y�p��/�����u뮺��[�J��Ǻ�U7�pUՊ�&��N���:r�s���5*F��)�\T6r���ff�ܡ�[',�����K闶#�۔��u ^{Q�OBXl�����D���Ƚwc	3pKo��X��n{0N�/�x>J��^��+/�V�ʕ�f֑����ξ��#��G���ohn*XS����� �����,\4�Q1� ���a�q�Y;v�og͚�0l�#F ��1c��,x\�4��𽧁�>g�k����A*����)������{��b�ͬ?Ʒk��Ҩ HM}<^;�X�.zf�������Nd�4^ح�+��ܰ�/x|�έa?��R=�&?�"kt��vw���<> �BM �K��<���9�X���͗�d����]5�X�����9Z�{O	�*.{�7>5{��򁱞�;w.2��w���2�L{�}ߑ�y{�̢��zpX8a36�1��R2c����������b$Q[7|�˥O������$��c����c�49������k9��FsCR�f\Ӥs4��⚌�ɵ�����":⡟]|�Xk�R�����o7b�Fٴ}��������54ԗ`ggӲx�B�c��cP()����P,����0�J�AJ�-��ƍ;�ZH�*���iih�k'l9I)���i����\*����-�3_������{���Z^���S�&ask�(���jb_H����4��$3vp~��^�#�v��?o���/�N7�ِ�$��Fk�Eẃuil�*��s}. �hѢ�ZH*cKaa���?#�|�ZJ�m����:s�����G�ϗ��� ��:5+��I8�;ƚ8ৱ�o[ǧ�=�~����?��=�s�wT�3mJ��LBDy�6Wr0j߮������)N�$#��?�?��|��kl{�$ca0^chw�N�b��eY�^={V�;|N(��y4�}�K�.��z=ƾ}�Vw���s�������s��Ds�����s�ҟ��O���K~�
ğ �C*.��{ܸZr�R�1R�H��k���%k*7L�������;�e*�����U�+V��éTH�j�y֑��{H�WY�X��x�IU�M��4_�.g�-uٶ�����ﭞ��b���c?[̧,��S��{�h��޿d�m��R)y޼yL�8�f�СG�U�r���\cg̘�^ "Rӽz�Z�E��"}z̏�}m�`-���y��iB����-��a�>=t`�[W����Ԡ��KW���s�[䤥�d�����.�]���Qip�Տ�.n{��b��UZ�ǎ̎C:���T�bѨ�Vr�g�ޫ��tK�9tC3M���VN|����H�r�/����k8J:H[.<��/�u�.<��ʝV�|c�a��i�J�xZE{ذa��f+��eYt���sJKK���k:uƒ9�}I�gn�,�ɆY���s�>;�_�Ѥ���t"��x�A���m��g��f��DS^2֨s.�=R6��􀑭��7k�I4K꒩"��Y�L�`_q陑.����Ā�S�<���JX5<�).fB�HI����Y����pF�ӻ�������q����3��,S_�z���i@屢�ֱŒ$%�ҏ~���V�j;��i��'�����W����|+��B��$���ϻ?:����7��Ly�XHS�����]�1�b݊fѺ �8��Fz`�^�v������_�lk�;���=Xcb�;�V��CZd�G�m��F[:�"�]}E[~�wPِ�C��p˸q;�ǭw�yg����/����0�G"��g�uֻ}��Y��Ͼ�aÆyMC&܋6��V�|s�S}��{����Z.�C��h�3�w:�׼KK�~�,^JNv�[�Bq3���Њ�[c^���Z���u�|��%�cI������(//'�K����������g��"�M�7�׌u�N^:�X��?B���G�c����?�2h�4o    IEND�B`�PK   6f�X����`  [  /   images/fc6d97d6-a1d8-4630-b4a2-8bef38b47130.png[��PNG

   IHDR   d   -   X���   	pHYs  �  ��iTS   tEXtSoftware www.inkscape.org��<  �IDATx��\tT��޼�QiԻ�PA	���b��[l��N�v�����ݜ�g�l��8�u�u�u��F�`0ŀ�$H �PA�޻FS���4B`p��q��#kt���������G\kN��G(�B?W�k�}�t��E?��s��n��ݕtnzw�Ӊ� _�d'@_�l6�t
4�C:����j��3�A&�D�G���1:j����^U�>00�Ŧ����胃�[AK���FY
��F1D?�*���0z�>2<*�p��󆇧F��Xen��^��2��Q�����d򄗷�|������t>>����6�S/�Ԑ��ޣ��@OϠד��9��p8�ݭ�=<��&���e�Fړ�c����tⁿ���p��uw�ႃ&���� f[��
���+Ve!vjm�7�������"19�5LQ`����ǽȞ33∩CB���/�����Db�F7�}���>���P�_�J�����8Dk1cɲLb��8}�{�DO��e6)�%��-����;s���L��;��:,�{�|����;8��$������E����L(�?��u�x���h^��"����X*N_�?<�T��t���G��Z<���$�`���7j�q��<��͢H$�.�a��2<���E�,l|CC�z� �
=k����XT8]�R�U��;����<u/MX��c;�����ˁ�����O֢�d=��@z��6�@ىP���w��l��w s�B�w��$����p��?@V&Y��'����?�BkK� 33]��:��/m|%zz��ޝ��e'K�{a݆�bm��BV����}{<p۝+�����F֌Q(d�����d1�ٹ3�Ghà1U�]���;�����CGkP0+g)V���[vczJ|�u�f -�&,_��m�� iZ7	O����,�=oݸ	S�I9T�1q���h�����jFp���B#���g�c���[��b�����&�0[6BϦ���CHN2`�r���l���>R�F1�[�ۉ�L�o��?ۈ��Q,]b�֭v��葖҅g�ڄ�(V��c�6;��TbP~��f���p��v��"g� ^x~1Ɓ���a�N;�U�����l#t`�Zv�&��̷���An��끽�2}`�";���"��7 )�y��eN��a�)x`��E
�8�z��w���,G���(U���Ě[Tlܼ�A�}�8S����Ik�Ӛ?�{�Z�u�*��������|�Z�~ˆ�V�F�À�
�u�	�u��,�@{s��ی�?r�9������wۈ'e�O#*z��-=�-��QzԞ���8\�Iww�#<��/�p����13����G�O46�PN��!����� �2<���*w�F]�9�HnjI��[��S4�F��x��o�}�F��9ȝ81/σ����J���R;��,X�'W7�AG�{#m�0�E��ޑ�`�E���;`A驯����%�mqa1������%7��Qb�i|_�--qS�JF���"e�ß�UW7Hn���q+������#(ȅ�3K�ﰢ���g�Qp�8�(Ą}����r�2��SPT��Q�e6z�AF� :Z'2��HƋ���I��S���1-AG�b�446��eV�[��ԩ:���b��4bz32�-X���)JAe�s榢�����p/����T[1sv2�dmx ����Y���H���G��^�|���E(Ng�н<��Y3�hvbl;��(@�Ҋ��hHoo)��+��|�0���&�0bq��6!HH���d��.Z�W�ɏ�v���
�5;0<b�=�^�p��z���L��D{N����[w�I�]��v�l��(�xU#�t�5-��={=p�Db|�x��d����z��,���Uথ�Pt$��\�<K�.2��(����B�;ɂH���13vG�

i"�78�m� FѠ)(�/B�4�՘�%Kc%�9\��SFH�p����'9r�bc����Ś��W&Y�q�#*�C�.�M%�>]�QQa��-!Xuk��s����b�U��X}k��x��|Z��)8]i���f�(.��*36J�(+��-krIV��XuAb�q�zM�쳕&��9B�:=�A�b��u�ƗxPM�C�Q���K(S!A�Q[[��rs�:,�9O�X���LW�ڮ�����ROMn�"{ɱs�U.̝�C�ω�D��҅g�܈Y��iI�h\|"�<��&AM�W�۱aJ��rc���M��Ĉٴ!;�iC�Cx��-��ƚ;�q�Ǭ�x#��_nAh�?�{��k�W�Y)�lv��y\b��~��w�oX nI�!N���;Bn�!�?^�g@h������"��)BOV2���ۋIH1��Y:�F����W�^^�LrA�y��P'���~y�&'Y���/DmM�y�$�Z����1`�T�_$2�I���"���'q�����G��#Y�#	�����8G�٠�^�A���n-�$�tٹ�ZhQF����B.�xB����TU6	]p6�y@FS/��-��3ol����thI��`�^NW����O����>��N����/���y�D0�j�W���
:�:��ʁ��*�F������in:���7���Wppfm|�p<�f:�s��ێ
_��e��g���*�;C��Ƈ�&�c.���pD���ϗ�3�ƫѵ���ҹ}S�;(����}���<�����O��J��``� ���$�2����� ��3�h.��?D��>��&4��T�×il9-ͽR�ȃq�	�նQ��C���s�;��c�RAA�$�
�܂��[����	C}J�|�T#��+j��왴Pܮhp���*�4�\m�XK��j1)���'�[#We���@.L�qU�M��a�P����{ ��dY������5)�8%�(R�c�tw_V��eQ������F�Ȍ��7�{0=-J\١��^��ukʗ0{e���+Ȅ�]�[���`�:�5���2s���\�|�e��6�]jY��{�����F�|Ė����u�(9�8
�a�f4����o���j��q	��zlf���Ȩ �,�X39�������' ��a�5��PO���BI��s(����ŗ\w��&(��gh��I9��Ж�+�'_wcXIa^*�b ��6tZ�P?}�l��+VgP��3)��{�`�����~��FF��8݄����t�mm*N�:��v���S�E ��E�1�U��ji�$�F�{1H��F�-�ɾx4����+lq�Ŋ>�S7ç�����J.��������4^��`�H����)��+qH}0!^��4��nL�L�Ŝ�dXH|���уw�*,}#�*����|�DV�e�p����a#sy�~蚖��1 ��ʤ�9`��lATL�d���
6!�`��5����~�=�u��������]��>o~2��%�X�a�$u
��Z���8���kb��YƵ�c����q��1����0�zbp@;�<[�,��O���'�l��w`��,-:	��?o@N^6���JyN��s�0�kAi����CMM1ҲnEP���1nD��<֤��q��G����>�V�F�#�>����ЖS	�>*y��,�m[�cf�}ؽ��,���!"�EG��������I|�ᒃ��tknU�8WQn<ALlv�v�Z�d+�J��zzE Z�� "Ҍ��~)G��<������[N�0V�� 2����`ܳ.[7���>��WV;�6]�Y�Td�Os��1z)�ݨM%���Q;`C���}*{�h�_�MOl,��P_DP���yTt A�.��iI�(o!q?J9���s��>�c�*gNbz�"e�y]lhGXd&}Q��+�$;�{�5E|�Z	�x����z���!�2ns�x����#�5���('֣c�k쫤�<�`pJO\�/�ir��.�#�?�PV\���X�c=����-�O�\���<�|I�?{j!~�ě��(��OȒ�Q����M#��v<�jF�� |���	����\��5z{���9(�⮻gS�݁��R�#n.9��D�I�?�H��CF���"`v�ArAY��������獦����w��ݷ����o����/v�0���o���}�P�N�iqJ��,apc�޷�B>��q�%.t���Y���(!쁯�l��,ET��]����U2�����Rp�8K�8Q^NҚ��ٳ%H�u	e9	)��;�Xrjv�Z���#������%�n:,Zg�~N�c��gYAYq���='�|p�7ٺ�O��~��G�ط��˹���1yj(��FY��ش�Nf�JJou�,;K��Z���
��Z��������[�
���q�sl��>�� �g��<=B��\�Mˈ�����N�%��ڱ%+�ʊ4��t-.�ݸm[�i(���u5LO�!+�PV���V¢�K(�k�\�5��o��ri�}�c�e<�gq���c��MÔ�`t�@8��%	� _�߯N2�=�	��(�(Cj���t�QY8SQ�U+U��0z�5UGYl�>�"����o��R�5�����/O^ aۻ�\�k~G� ��;��d9u�(<24*�^.8�hJM(+��/$2ʊ�U0u�(k��b��w>2�o%�gAX�i��?���H\P�͆��
�|�(?o��ߴ�k`�����n�ģg��_��x����P���U�&e����f��<PI(���F$��0�QV����z��)��ЁN�t��]`��B��F!��
-����5�cTyv��K�^�{��|���V<�ʮv �e�]c7�9��-�Ύ>x�gQ�(�P�A���PR\��,��Z�6+��yP
��p@��n����~w�݇��/rNM�0��t�&}��wSFpi�N	�«���F����iBY?�QŐrs�����P��q���E��)fn��E=��1w?	��.TW�~D
�gL^��X��̘?c(�T�E���O|���'��c�҄��#˰ck�/!�PVcC�g.vl+�g����%G�0=5J&��ű��,�}_KK���P�Oe8.x{e�eDPy��i�t��y�`�*���X�ͦs��;Vܬ�Ty)Rg,�tb�i��z$�Z��"�0˵��Zy��4|Di�:���O|��nv�ki�>r����?Kʆ�
�3���.��_�(zP�I��K9F��`m1ʊ������	eM���>Ϥ�x�!~�L��XS(P]�>��7c}l$(o��Y�c1^��5�g#�jW9�1d�]�dE��3g��Ȳu�8<�K�x��$�s��<d��K �Ok|�v�Bv�*�[$�iQr�s��`RX��h��q�`0x�l��W	�*�����K���>�@�̾Z��h��c�L]XP+&x�=���.ŷ=���_�~�!��{���EPo�v�}{�����f1bb)s�sߺ�8�Y?Gn�-:'���戀6�w���I���娮n%�D��_��r1��3Υ�z�H��׻��
�`���*Q���2������ʻ��CH�/0u��HH�+,.�����z.��2��r�����gD�gv-4�,����b��9 �3rc���p0d7x����BZt�V�>vJ~�����_��S���K�x�tdω���G��=8v�Ԓ2=B��?��[�WU�q�j��"?�}R�O�{�Ճr+>9m�(p�|#�W!�`�\�����{�6*_�fjw���)'����1k>C`�^p�
K���Ƹ���*sf� v�|I\'�E�~�ң��ʡ���B���Yj\B�N\��n^N�)c���o��p��t�'o�_�IY˙In+`�)��9(�z[�\YMI��L�3]�3�ٍ�X�!��B�g�FU��}ߙ'�ow��f�s#w�y��;�\�௷)�Wu���e7R��@��Ä���H��/{��F��|�\ǃ����QԒ�b��G�܁��kq�9<��	�o�V�[�d���q���T�����eS��*���Gq�������$7��������$��=Xʧ��*��������_��^��@�G:;�v=��,�\-u_*���DmM�\������>�����&qU|]S�����8�✉����EP�δ���v}-D� 2g����o>p�O�E�Wܾ���m!���3?�Մ)ɰ��x�t��K�k9�X馃��D��G�Lg�r��Mh_IQ'���&~��W~�������.+ٸ��w���y�E#��C    IEND�B`�PK   6f�Xږ�5[  �(     jsons/user_defined.json�Z�n�H�AO=���}ɛm3F;Kۙ���jcB�L��$H���$�8qQ)�i�`X"�ܪ�=�ι�����2N_L���bQV1Lg��q�.\��|�޺�������?���؋Uؖ�b���/�&�7/'w�Z��m�La����q��
c���@�|�~6- f�4F!�0F<F���E���^G'l��xX.�Xm��Gg���x/6�m�1�<���\nڅ<��m�᳧Apl0�E �{O!�
�j���G,�e�ƕ~Q���*�fܠc�8�E(�a��$���`?ƛ���?�?����"\]��uU,�/�M��C^��s��j1_׻�2E��p���ŗ��ʰ������V�_[XTu�6���S�oX��:��r^�
�1-��IM3b�����E�?-V0z�ys�b=`�}֍Mlz���up�����Y���	�\$�r<p�����U���	�ܤ�㡓���ho�������)K�x�)K�x�)K�x�)K�x�)K�x�)K�x�)K�x�)K�hഃ�x<����Q�r��GR�����R��u M�JFT4�*QД�d�
IS���J$�8TϨ����}�Z�/�
��w�j�X�զlL�}=�_}��2����-��3���mBcIT0Ð3^ �F�q�S�&�b橥`����$
q�26z�"����8���ϖ��v��nj3�٭�'�pR�7v�y���fxftN����b݄�7���� �B�:���#2N�0Ǧ�x��<��mr"uR83�@��23����J����c�L?y>�-C�>�9��A:��SXʂ3���������z��̡�ÇeU[l;����m	�q�s��_�TW�u��΋�庬��n��6��<��Q
g�ma�f�j�~�"�b�-7��*l�10��O�˥��n8e�?P����c�-�
�8�YZX�QNN��7��ǯ*$�K�Á"M��B���6���❅�F�L�G��r���L+�iW�� ��S{X� �`&�bppA� �r�0��~@瀝D������P��̀��~��ܣ+��;D{Q"�
Jҡp�k8�4�5C��N����R� ��H���V"�"�2Y��\��p�sf,�՛q��~#��%�P��gS�g�y��ŕ<��&2�V3a2l@�gı���1|�i�^���N�j�/I/��WW�f��U>�m��7"' �Aڧ�hCu��ȉ��*E��9��Pm����앩[8�� �!.�E�Qg9��p���Y~$���M����B�l}��bDg`^�Fi��ǜ(�wwR����Rz���χ�[�cO)�r8���J=��A��3�i��/�倶�>��h�<|��a���5�9�&.='�����$��=������%g�9��C��F�jH{��A���iG���A��{��}�&�W��Q"B=Y�(�"�k
���q�cp�	�����|�ys��HL'��W�E�ƪhXO&�̣�1�	h��Qо"�*�"	)��D��EBY2��TIj9]x�
�M� �F��Z�ǂi�ayZ��	&x�bV׸�U�Jf
��qP�Tr|�E��-��<c5>��W:�j{���f̨���U��> u ��)3ywu3@ڰ�Ig��?���p%O� m�� ��U��}��S�7����x�Հ���4������ܜ��#��C��\����1U�)g���?�aU�%fh�G������)��������1��g��ʎ�$iS��O����L�ۦ���������oK`���=�:�V���6V/�M�1՟c��$�-�T��]U�k��R�gLk`����o^����R��@wN�ū#\��,�#���PK
   6f�Xn�
�$  ��                  cirkitFile.jsonPK
   6f�XG�~��  � /             �$  images/0739a1b1-a163-452a-a325-ab452d55b136.pngPK
   6f�X�;�К> � /             ��  images/277be1dd-7489-4b2a-8eff-ec6391927629.pngPK
   ,V�X&�n�-u  #u  /             �$ images/294439aa-ec9f-4672-895d-838110657847.pngPK
   6f�X�j�� 7q /             � images/3afa6c98-60d7-4a37-9aec-be07fd386e0e.pngPK
   V�X.D��N �M /             z
 images/4f771273-f62d-49a2-b0d2-ce9da7065853.pngPK
   ,V�X:�I��  �  /             �� images/65cd5dc4-66ed-44a6-97e2-8bf96ed14d67.pngPK
   vb�X��n} � /             "[ images/87fd8349-f00c-446b-9712-cb30a7c611c5.pngPK
   6f�X	�\  \  /             q� images/898ac7d1-13d0-4a1b-8b5c-ab7066f4327a.pngPK
   6f�X�Ƚ׌  �  /             � images/9185dcb2-65ea-4de0-8d42-42cedb1b5634.pngPK
   vb�XT�7Pb #y /             �� images/c2d54090-2fd1-4cc2-9c7d-28b872c3ce05.pngPK
   V�X+���q6 X6 /             �` images/d8919090-1cba-41eb-9d62-14d110867e7b.pngPK
   6f�X����`  [  /             N� images/fc6d97d6-a1d8-4630-b4a2-8bef38b47130.pngPK
   6f�Xږ�5[  �(               �� jsons/user_defined.jsonPK      �  ��   